//
// Verilog description for cell floating_point_multiplication, 
// Thu Dec 12 13:40:37 2019
//
// LeonardoSpectrum Level 3, 2009a.6 
//


module floating_point_multiplication ( input_a, input_b, product, underflow, 
                                       overflow ) ;

    input [31:0]input_a ;
    input [31:0]input_b ;
    output [31:0]product ;
    output underflow ;
    output overflow ;

    wire nx12, nx26, nx42, nx56, nx74, nx88, nx104, nx118, nx138, nx152, nx168, 
         nx182, nx200, nx214, nx230, nx244, nx252, nx290, nx292, nx322, nx326, 
         nx362, nx364, nx418, nx422, nx490, nx492, nx570, nx574, nx674, nx676, 
         nx778, nx782, nx914, nx916, nx1042, nx1046, nx1210, nx1212, nx1362, 
         nx1366, nx1562, nx1564, nx1738, nx1742, nx1970, nx1972, nx2170, nx2174, 
         nx2434, nx2436, nx2658, nx2662, nx2954, nx2956, nx3190, nx3192, nx3208, 
         nx3212, nx3214, nx3218, nx3220, nx3224, nx3226, nx3230, nx3232, nx3236, 
         nx3238, nx3242, nx3244, nx3248, nx3250, nx3254, nx3256, nx3260, nx3262, 
         nx3266, nx3268, nx3272, nx3274, nx3278, nx3280, nx3284, nx3286, nx3290, 
         nx3292, nx3296, nx3298, nx3302, nx3304, nx3308, nx3310, nx3314, nx3316, 
         nx3320, nx3322, nx3324, nx3530, nx3532, nx3796, nx3800, nx3804, nx3806, 
         nx3810, nx3812, nx3816, nx3818, nx3822, nx3824, nx3828, nx3830, nx3834, 
         nx3836, nx3840, nx3842, nx3846, nx3848, nx3852, nx3854, nx3858, nx3860, 
         nx3864, nx3866, nx3870, nx3872, nx3876, nx3878, nx3882, nx3884, nx3888, 
         nx3890, nx3894, nx3896, nx3900, nx3902, nx3906, nx3908, nx3912, nx3914, 
         nx3918, nx3920, nx3928, nx3946, nx3968, nx3992, nx4010, nx4014, nx4020, 
         nx4030, nx4038, nx4046, nx4054, nx4062, nx4070, nx4078, nx4086, nx4094, 
         nx4102, nx4110, nx4118, nx4126, nx4134, nx4142, nx4150, nx4158, nx4166, 
         nx4174, nx4182, nx4190, nx4202, nx4210, nx4218, nx4226, nx4234, nx4242, 
         nx4250, nx4258, nx4266, nx4274, nx4288, nx4290, nx4294, nx4302, nx4304, 
         nx4322, nx4324, nx4342, nx4344, nx4362, nx4364, nx4382, nx4384, nx4402, 
         nx4404, nx4422, nx4424, nx4442, nx4444, nx4462, nx4464, nx4482, nx4484, 
         nx4590, nx4592, nx4598, nx4600, nx4620, nx4622, nx4640, nx4642, nx4660, 
         nx4662, nx4680, nx4682, nx4700, nx4702, nx4720, nx4722, nx4740, nx4742, 
         nx4760, nx4762, nx4780, nx4782, nx4884, nx4896, nx4904, nx4906, nx4924, 
         nx4926, nx4944, nx4946, nx4964, nx4966, nx4984, nx4986, nx5004, nx5006, 
         nx5024, nx5026, nx5044, nx5046, nx5064, nx5066, nx5164, nx5166, nx5172, 
         nx5174, nx5194, nx5196, nx5214, nx5216, nx5234, nx5236, nx5254, nx5256, 
         nx5274, nx5276, nx5294, nx5296, nx5314, nx5316, nx5334, nx5336, nx5430, 
         nx5442, nx5450, nx5452, nx5470, nx5472, nx5490, nx5492, nx5510, nx5512, 
         nx5530, nx5532, nx5550, nx5552, nx5570, nx5572, nx5590, nx5592, nx5682, 
         nx5684, nx5690, nx5692, nx5712, nx5714, nx5732, nx5734, nx5752, nx5754, 
         nx5772, nx5774, nx5792, nx5794, nx5812, nx5814, nx5832, nx5834, nx5920, 
         nx5928, nx5932, nx5940, nx5942, nx5960, nx5962, nx5980, nx5982, nx6000, 
         nx6002, nx6020, nx6022, nx6040, nx6042, nx6060, nx6062, nx6144, nx6146, 
         nx6152, nx6154, nx6174, nx6176, nx6194, nx6196, nx6214, nx6216, nx6234, 
         nx6236, nx6254, nx6256, nx6274, nx6276, nx6354, nx6366, nx6374, nx6376, 
         nx6394, nx6396, nx6414, nx6416, nx6434, nx6436, nx6454, nx6456, nx6474, 
         nx6476, nx6550, nx6552, nx6558, nx6560, nx6580, nx6582, nx6600, nx6602, 
         nx6620, nx6622, nx6640, nx6642, nx6660, nx6662, nx6732, nx6744, nx6752, 
         nx6754, nx6772, nx6774, nx6792, nx6794, nx6812, nx6814, nx6832, nx6834, 
         nx6900, nx6902, nx6908, nx6910, nx6930, nx6932, nx6950, nx6952, nx6970, 
         nx6972, nx6990, nx6992, nx7054, nx7062, nx7066, nx7074, nx7076, nx7094, 
         nx7096, nx7114, nx7116, nx7134, nx7136, nx7194, nx7196, nx7202, nx7204, 
         nx7224, nx7226, nx7244, nx7246, nx7264, nx7266, nx7320, nx7332, nx7340, 
         nx7342, nx7360, nx7362, nx7380, nx7382, nx7432, nx7434, nx7440, nx7442, 
         nx7462, nx7464, nx7482, nx7484, nx7530, nx7542, nx7550, nx7552, nx7570, 
         nx7572, nx7614, nx7616, nx7622, nx7624, nx7644, nx7646, nx7684, nx7692, 
         nx7696, nx7704, nx7706, nx7740, nx7742, nx7748, nx7750, nx7782, nx7794, 
         nx7810, nx7812, nx7824, nx7826, nx7832, nx7836, nx7840, nx7844, nx7856, 
         nx7860, nx7864, nx7868, nx7880, nx7884, nx7888, nx7892, nx7904, nx7908, 
         nx7912, nx7920, nx7926, nx7932, nx7938, nx7944, nx7950, nx7956, nx7962, 
         nx7970, nx7974, nx7976, nx7980, nx7982, nx7986, nx7988, nx7992, nx7994, 
         nx7998, nx8000, nx8004, nx8006, nx8010, nx8012, nx8016, nx8028, nx8040, 
         nx8048, nx8054, nx8066, nx8074, nx8080, nx8092, nx8100, nx8106, nx8136, 
         nx8142, nx8144, nx8150, nx8158, nx8170, nx8178, nx8184, nx8214, nx8220, 
         nx8222, nx8228, nx8236, nx8248, nx8256, nx8262, nx8292, nx8298, nx8300, 
         nx8306, nx8314, nx8326, nx8334, nx8340, nx8370, nx8376, nx8378, nx8384, 
         nx8392, nx8404, nx8412, nx8418, nx8448, nx8454, nx8456, nx8462, nx8470, 
         nx8482, nx8490, nx8496, nx8526, nx8532, nx8534, nx8540, nx8548, nx8560, 
         nx8568, nx8574, nx8598, nx8604, nx8610, nx8614, nx8620, nx8624, nx8638, 
         nx8652, nx8666, nx8680, nx8694, nx8714, nx8720, nx8726, nx8732, nx8738, 
         nx8746, nx8750, nx8754, nx8776, nx8794, nx8812, nx8842, nx8848, nx8878, 
         nx8884, nx1245, nx1247, nx1251, nx1253, nx1255, nx1257, nx1259, nx1261, 
         nx1265, nx1267, nx1269, nx1271, nx1273, nx1275, nx1277, nx1279, nx1281, 
         nx1285, nx1289, nx1293, nx1299, nx1301, nx1303, nx1305, nx1307, nx1309, 
         nx1311, nx1317, nx1323, nx1329, nx1331, nx1333, nx1335, nx1341, nx1343, 
         nx1349, nx1359, nx1367, nx1375, nx1383, nx1391, nx1399, nx1407, nx1415, 
         nx1423, nx1431, nx1433, nx1435, nx1441, nx1445, nx1449, nx1453, nx1457, 
         nx1461, nx1465, nx1469, nx1473, nx1477, nx1481, nx1485, nx1489, nx1493, 
         nx1497, nx1501, nx1505, nx1509, nx1513, nx1517, nx1519, nx1525, nx1527, 
         nx1529, nx1531, nx1533, nx1535, nx1537, nx1539, nx1541, nx1543, nx1545, 
         nx1547, nx1549, nx1551, nx1553, nx1555, nx1557, nx1559, nx1561, nx1563, 
         nx1565, nx1567, nx1569, nx1571, nx1573, nx1575, nx1577, nx1579, nx1581, 
         nx1583, nx1585, nx1587, nx1589, nx1591, nx1593, nx1595, nx1601, nx1609, 
         nx1611, nx1613, nx1615, nx1617, nx1619, nx1621, nx1623, nx1625, nx1629, 
         nx1631, nx1635, nx1641, nx1649, nx1651, nx1653, nx1655, nx1657, nx1659, 
         nx1661, nx1663, nx1669, nx1677, nx1679, nx1681, nx1683, nx1685, nx1687, 
         nx1689, nx1691, nx1697, nx1705, nx1707, nx1709, nx1711, nx1713, nx1715, 
         nx1717, nx1719, nx1725, nx1733, nx1735, nx1737, nx1739, nx1741, nx1743, 
         nx1745, nx1747, nx1753, nx1761, nx1763, nx1765, nx1767, nx1769, nx1771, 
         nx1773, nx1775, nx1781, nx1789, nx1791, nx1793, nx1795, nx1797, nx1799, 
         nx1801, nx1803, nx1809, nx1817, nx1819, nx1821, nx1823, nx1825, nx1827, 
         nx1829, nx1831, nx1837, nx1845, nx1847, nx1849, nx1851, nx1853, nx1855, 
         nx1857, nx1859, nx1865, nx1873, nx1875, nx1877, nx1879, nx1881, nx1883, 
         nx1885, nx1887, nx1889, nx1893, nx1901, nx1903, nx1905, nx1907, nx1909, 
         nx1911, nx1913, nx1915, nx1917, nx1919, nx1921, nx1923, nx1925, nx1927, 
         nx1929, nx1931, nx1933, nx1935, nx1937, nx1939, nx1941, nx1943, nx1945, 
         nx1947, nx1949, nx1951, nx1953, nx1955, nx1957, nx1959, nx1961, nx1963, 
         nx1965, nx1967, nx1969, nx1971, nx1973, nx1981, nx1983, nx1985, nx1987, 
         nx1989, nx1991, nx1999, nx2001, nx2007, nx2009, nx2015, nx2021, nx2027, 
         nx2029, nx2031, nx2033, nx2035, nx2037, nx2039, nx2041, nx2047, nx2053, 
         nx2055, nx2057, nx2059, nx2061, nx2063, nx2065, nx2067, nx2073, nx2079, 
         nx2081, nx2083, nx2085, nx2087, nx2089, nx2091, nx2093, nx2099, nx2105, 
         nx2107, nx2109, nx2111, nx2113, nx2115, nx2117, nx2119, nx2125, nx2131, 
         nx2133, nx2135, nx2137, nx2139, nx2141, nx2143, nx2145, nx2151, nx2157, 
         nx2159, nx2161, nx2163, nx2165, nx2167, nx2169, nx2171, nx2177, nx2183, 
         nx2185, nx2187, nx2189, nx2191, nx2193, nx2195, nx2197, nx2203, nx2209, 
         nx2211, nx2213, nx2215, nx2217, nx2219, nx2221, nx2223, nx2229, nx2235, 
         nx2237, nx2239, nx2241, nx2243, nx2245, nx2247, nx2249, nx2251, nx2255, 
         nx2261, nx2263, nx2269, nx2271, nx2273, nx2275, nx2277, nx2279, nx2281, 
         nx2283, nx2285, nx2287, nx2289, nx2291, nx2293, nx2295, nx2297, nx2299, 
         nx2301, nx2303, nx2305, nx2307, nx2309, nx2311, nx2313, nx2315, nx2317, 
         nx2319, nx2321, nx2323, nx2325, nx2327, nx2329, nx2331, nx2339, nx2341, 
         nx2343, nx2345, nx2347, nx2349, nx2357, nx2359, nx2361, nx2363, nx2365, 
         nx2367, nx2369, nx2371, nx2373, nx2375, nx2377, nx2379, nx2381, nx2383, 
         nx2385, nx2387, nx2389, nx2395, nx2401, nx2407, nx2413, nx2415, nx2417, 
         nx2419, nx2421, nx2423, nx2425, nx2427, nx2433, nx2439, nx2441, nx2443, 
         nx2445, nx2447, nx2449, nx2451, nx2453, nx2459, nx2465, nx2467, nx2469, 
         nx2471, nx2473, nx2475, nx2477, nx2479, nx2485, nx2491, nx2493, nx2495, 
         nx2497, nx2499, nx2501, nx2503, nx2505, nx2511, nx2517, nx2519, nx2521, 
         nx2523, nx2525, nx2527, nx2529, nx2531, nx2537, nx2543, nx2545, nx2547, 
         nx2549, nx2551, nx2553, nx2555, nx2557, nx2563, nx2569, nx2571, nx2573, 
         nx2575, nx2577, nx2579, nx2581, nx2583, nx2589, nx2595, nx2597, nx2599, 
         nx2601, nx2603, nx2605, nx2607, nx2609, nx2611, nx2615, nx2621, nx2627, 
         nx2629, nx2631, nx2633, nx2635, nx2637, nx2639, nx2641, nx2643, nx2645, 
         nx2647, nx2649, nx2651, nx2653, nx2655, nx2657, nx2659, nx2661, nx2663, 
         nx2665, nx2667, nx2669, nx2671, nx2673, nx2675, nx2677, nx2679, nx2681, 
         nx2683, nx2685, nx2687, nx2689, nx2697, nx2699, nx2701, nx2703, nx2705, 
         nx2707, nx2715, nx2717, nx2719, nx2721, nx2723, nx2725, nx2727, nx2729, 
         nx2731, nx2733, nx2735, nx2737, nx2739, nx2741, nx2743, nx2745, nx2747, 
         nx2749, nx2751, nx2753, nx2755, nx2757, nx2759, nx2761, nx2763, nx2765, 
         nx2767, nx2769, nx2771, nx2773, nx2775, nx2781, nx2787, nx2793, nx2799, 
         nx2801, nx2803, nx2805, nx2807, nx2809, nx2811, nx2813, nx2819, nx2825, 
         nx2827, nx2829, nx2831, nx2833, nx2835, nx2837, nx2839, nx2845, nx2851, 
         nx2853, nx2855, nx2857, nx2859, nx2861, nx2863, nx2865, nx2871, nx2877, 
         nx2879, nx2881, nx2883, nx2885, nx2887, nx2889, nx2891, nx2897, nx2903, 
         nx2905, nx2907, nx2909, nx2911, nx2913, nx2915, nx2917, nx2923, nx2929, 
         nx2931, nx2933, nx2935, nx2937, nx2939, nx2941, nx2943, nx2949, nx2955, 
         nx2957, nx2959, nx2961, nx2963, nx2965, nx2967, nx2969, nx2971, nx2975, 
         nx2981, nx2983, nx2985, nx2987, nx2989, nx2991, nx2993, nx2995, nx2997, 
         nx2999, nx3001, nx3003, nx3005, nx3007, nx3009, nx3011, nx3013, nx3015, 
         nx3017, nx3019, nx3021, nx3023, nx3025, nx3027, nx3029, nx3031, nx3033, 
         nx3035, nx3037, nx3039, nx3041, nx3043, nx3045, nx3047, nx3055, nx3057, 
         nx3059, nx3061, nx3063, nx3065, nx3073, nx3075, nx3077, nx3079, nx3081, 
         nx3083, nx3085, nx3087, nx3089, nx3091, nx3093, nx3095, nx3097, nx3099, 
         nx3101, nx3103, nx3105, nx3107, nx3109, nx3111, nx3113, nx3115, nx3117, 
         nx3119, nx3121, nx3123, nx3125, nx3127, nx3129, nx3131, nx3133, nx3135, 
         nx3137, nx3139, nx3141, nx3143, nx3145, nx3147, nx3149, nx3151, nx3153, 
         nx3155, nx3157, nx3159, nx3161, nx3167, nx3173, nx3179, nx3185, nx3187, 
         nx3189, nx3191, nx3193, nx3195, nx3197, nx3199, nx3205, nx3211, nx3213, 
         nx3215, nx3217, nx3219, nx3221, nx3223, nx3225, nx3231, nx3237, nx3239, 
         nx3241, nx3243, nx3245, nx3247, nx3249, nx3251, nx3257, nx3263, nx3265, 
         nx3267, nx3269, nx3271, nx3273, nx3275, nx3277, nx3283, nx3289, nx3291, 
         nx3293, nx3295, nx3297, nx3299, nx3301, nx3303, nx3309, nx3315, nx3317, 
         nx3319, nx3321, nx3323, nx3325, nx3327, nx3329, nx3331, nx3335, nx3341, 
         nx3343, nx3349, nx3351, nx3353, nx3355, nx3357, nx3359, nx3361, nx3363, 
         nx3365, nx3367, nx3369, nx3371, nx3373, nx3375, nx3377, nx3379, nx3381, 
         nx3383, nx3385, nx3387, nx3389, nx3391, nx3393, nx3395, nx3397, nx3399, 
         nx3401, nx3403, nx3405, nx3413, nx3415, nx3417, nx3419, nx3421, nx3423, 
         nx3431, nx3433, nx3435, nx3437, nx3439, nx3441, nx3443, nx3445, nx3447, 
         nx3449, nx3451, nx3453, nx3455, nx3457, nx3459, nx3461, nx3463, nx3465, 
         nx3467, nx3469, nx3471, nx3473, nx3475, nx3477, nx3479, nx3481, nx3483, 
         nx3485, nx3487, nx3489, nx3491, nx3493, nx3495, nx3497, nx3499, nx3501, 
         nx3503, nx3505, nx3507, nx3509, nx3511, nx3513, nx3515, nx3517, nx3519, 
         nx3521, nx3523, nx3525, nx3527, nx3529, nx3531, nx3533, nx3535, nx3537, 
         nx3539, nx3541, nx3543, nx3545, nx3547, nx3553, nx3559, nx3565, nx3571, 
         nx3573, nx3575, nx3577, nx3579, nx3581, nx3583, nx3585, nx3591, nx3597, 
         nx3599, nx3601, nx3603, nx3605, nx3607, nx3609, nx3611, nx3617, nx3623, 
         nx3625, nx3627, nx3629, nx3631, nx3633, nx3635, nx3637, nx3643, nx3649, 
         nx3651, nx3653, nx3655, nx3657, nx3659, nx3661, nx3663, nx3669, nx3675, 
         nx3677, nx3679, nx3681, nx3683, nx3685, nx3687, nx3689, nx3691, nx3695, 
         nx3701, nx3707, nx3709, nx3711, nx3713, nx3715, nx3717, nx3719, nx3721, 
         nx3723, nx3725, nx3727, nx3729, nx3731, nx3733, nx3735, nx3737, nx3739, 
         nx3741, nx3743, nx3745, nx3747, nx3749, nx3751, nx3753, nx3755, nx3757, 
         nx3759, nx3761, nx3763, nx3771, nx3773, nx3775, nx3777, nx3779, nx3781, 
         nx3789, nx3791, nx3793, nx3795, nx3797, nx3799, nx3801, nx3803, nx3805, 
         nx3807, nx3809, nx3811, nx3813, nx3815, nx3817, nx3819, nx3821, nx3823, 
         nx3825, nx3827, nx3829, nx3831, nx3833, nx3835, nx3837, nx3839, nx3841, 
         nx3843, nx3845, nx3847, nx3849, nx3851, nx3853, nx3855, nx3857, nx3859, 
         nx3861, nx3863, nx3865, nx3867, nx3869, nx3871, nx3873, nx3875, nx3877, 
         nx3879, nx3881, nx3883, nx3885, nx3887, nx3889, nx3891, nx3893, nx3895, 
         nx3897, nx3899, nx3901, nx3903, nx3905, nx3907, nx3909, nx3911, nx3913, 
         nx3915, nx3917, nx3919, nx3921, nx3923, nx3925, nx3927, nx3929, nx3931, 
         nx3933, nx3939, nx3945, nx3951, nx3957, nx3959, nx3961, nx3963, nx3965, 
         nx3967, nx3969, nx3971, nx3977, nx3983, nx3985, nx3987, nx3989, nx3991, 
         nx3993, nx3995, nx3997, nx4003, nx4009, nx4011, nx4013, nx4015, nx4017, 
         nx4019, nx4021, nx4023, nx4029, nx4035, nx4037, nx4039, nx4041, nx4043, 
         nx4045, nx4047, nx4049, nx4051, nx4055, nx4061, nx4063, nx4065, nx4067, 
         nx4069, nx4071, nx4073, nx4075, nx4077, nx4079, nx4081, nx4083, nx4085, 
         nx4087, nx4089, nx4091, nx4093, nx4095, nx4097, nx4099, nx4101, nx4103, 
         nx4105, nx4107, nx4109, nx4111, nx4113, nx4115, nx4117, nx4119, nx4121, 
         nx4129, nx4131, nx4133, nx4135, nx4137, nx4139, nx4147, nx4149, nx4151, 
         nx4153, nx4155, nx4157, nx4159, nx4161, nx4163, nx4165, nx4167, nx4169, 
         nx4171, nx4173, nx4175, nx4177, nx4179, nx4181, nx4183, nx4185, nx4187, 
         nx4189, nx4191, nx4193, nx4195, nx4197, nx4199, nx4201, nx4203, nx4205, 
         nx4207, nx4209, nx4211, nx4213, nx4215, nx4217, nx4219, nx4221, nx4223, 
         nx4225, nx4227, nx4229, nx4231, nx4233, nx4235, nx4237, nx4239, nx4241, 
         nx4243, nx4245, nx4247, nx4249, nx4251, nx4253, nx4255, nx4257, nx4259, 
         nx4261, nx4263, nx4265, nx4267, nx4269, nx4271, nx4273, nx4275, nx4277, 
         nx4279, nx4281, nx4283, nx4285, nx4287, nx4289, nx4291, nx4293, nx4295, 
         nx4297, nx4299, nx4301, nx4303, nx4305, nx4307, nx4309, nx4311, nx4313, 
         nx4315, nx4317, nx4319, nx4325, nx4331, nx4337, nx4343, nx4345, nx4347, 
         nx4349, nx4351, nx4353, nx4355, nx4357, nx4363, nx4369, nx4371, nx4373, 
         nx4375, nx4377, nx4379, nx4381, nx4383, nx4389, nx4395, nx4397, nx4399, 
         nx4401, nx4403, nx4405, nx4407, nx4409, nx4411, nx4415, nx4421, nx4423, 
         nx4429, nx4431, nx4433, nx4435, nx4437, nx4439, nx4441, nx4443, nx4445, 
         nx4447, nx4449, nx4451, nx4453, nx4455, nx4457, nx4459, nx4461, nx4463, 
         nx4465, nx4467, nx4469, nx4471, nx4473, nx4475, nx4477, nx4479, nx4487, 
         nx4489, nx4491, nx4493, nx4495, nx4497, nx4505, nx4507, nx4509, nx4511, 
         nx4513, nx4515, nx4517, nx4519, nx4521, nx4523, nx4525, nx4527, nx4529, 
         nx4531, nx4533, nx4535, nx4537, nx4539, nx4541, nx4543, nx4545, nx4547, 
         nx4549, nx4551, nx4553, nx4555, nx4557, nx4559, nx4561, nx4563, nx4565, 
         nx4567, nx4569, nx4571, nx4573, nx4575, nx4577, nx4579, nx4581, nx4583, 
         nx4585, nx4587, nx4589, nx4591, nx4593, nx4595, nx4597, nx4599, nx4601, 
         nx4603, nx4605, nx4607, nx4609, nx4611, nx4613, nx4615, nx4617, nx4619, 
         nx4621, nx4623, nx4625, nx4627, nx4629, nx4631, nx4633, nx4635, nx4637, 
         nx4639, nx4641, nx4643, nx4645, nx4647, nx4649, nx4651, nx4653, nx4655, 
         nx4657, nx4659, nx4661, nx4663, nx4665, nx4667, nx4669, nx4671, nx4673, 
         nx4675, nx4677, nx4679, nx4681, nx4683, nx4685, nx4687, nx4689, nx4691, 
         nx4693, nx4695, nx4697, nx4699, nx4701, nx4703, nx4705, nx4711, nx4717, 
         nx4723, nx4729, nx4731, nx4733, nx4735, nx4737, nx4739, nx4741, nx4743, 
         nx4749, nx4755, nx4757, nx4759, nx4761, nx4763, nx4765, nx4767, nx4769, 
         nx4771, nx4775, nx4781, nx4787, nx4789, nx4791, nx4793, nx4795, nx4797, 
         nx4799, nx4801, nx4803, nx4805, nx4807, nx4809, nx4811, nx4813, nx4815, 
         nx4817, nx4819, nx4821, nx4823, nx4825, nx4827, nx4829, nx4831, nx4833, 
         nx4835, nx4837, nx4845, nx4847, nx4849, nx4851, nx4853, nx4855, nx4863, 
         nx4865, nx4867, nx4869, nx4871, nx4873, nx4875, nx4877, nx4879, nx4881, 
         nx4883, nx4885, nx4887, nx4889, nx4891, nx4893, nx4895, nx4897, nx4899, 
         nx4901, nx4903, nx4905, nx4907, nx4909, nx4911, nx4913, nx4915, nx4917, 
         nx4919, nx4921, nx4923, nx4925, nx4927, nx4929, nx4931, nx4933, nx4935, 
         nx4937, nx4939, nx4941, nx4943, nx4945, nx4947, nx4949, nx4951, nx4953, 
         nx4955, nx4957, nx4959, nx4961, nx4963, nx4965, nx4967, nx4969, nx4971, 
         nx4973, nx4975, nx4977, nx4979, nx4981, nx4983, nx4985, nx4987, nx4989, 
         nx4991, nx4993, nx4995, nx4997, nx4999, nx5001, nx5003, nx5005, nx5007, 
         nx5009, nx5011, nx5013, nx5015, nx5017, nx5019, nx5021, nx5023, nx5025, 
         nx5027, nx5029, nx5031, nx5033, nx5035, nx5037, nx5039, nx5041, nx5043, 
         nx5045, nx5047, nx5049, nx5051, nx5053, nx5055, nx5057, nx5059, nx5061, 
         nx5063, nx5065, nx5067, nx5069, nx5071, nx5073, nx5075, nx5077, nx5079, 
         nx5081, nx5083, nx5085, nx5087, nx5089, nx5091, nx5097, nx5103, nx5109, 
         nx5115, nx5117, nx5119, nx5121, nx5123, nx5125, nx5127, nx5129, nx5131, 
         nx5135, nx5141, nx5143, nx5147, nx5149, nx5151, nx5153, nx5155, nx5157, 
         nx5159, nx5161, nx5163, nx5165, nx5167, nx5169, nx5171, nx5173, nx5175, 
         nx5177, nx5179, nx5181, nx5183, nx5185, nx5187, nx5189, nx5191, nx5193, 
         nx5201, nx5203, nx5205, nx5207, nx5209, nx5211, nx5213, nx5215, nx5217, 
         nx5219, nx5221, nx5223, nx5225, nx5227, nx5229, nx5231, nx5233, nx5235, 
         nx5237, nx5239, nx5241, nx5243, nx5245, nx5247, nx5249, nx5251, nx5253, 
         nx5255, nx5257, nx5259, nx5261, nx5263, nx5265, nx5267, nx5269, nx5271, 
         nx5273, nx5275, nx5277, nx5279, nx5281, nx5283, nx5285, nx5287, nx5289, 
         nx5291, nx5293, nx5295, nx5297, nx5299, nx5301, nx5303, nx5305, nx5307, 
         nx5309, nx5311, nx5321, nx5323, nx5325, nx5327, nx5329, nx5331, nx5333, 
         nx5335, nx5337, nx5339, nx5341, nx5343, nx5345, nx5347, nx5349, nx5351, 
         nx5353, nx5355, nx5357, nx5359, nx5361, nx5363, nx5365, nx5367, nx5369, 
         nx5371, nx5379, nx5381, nx5383, nx5385, nx5387, nx5389, nx5391, nx5393, 
         nx5395, nx5397, nx5399, nx5401, nx5403, nx5405, nx5407, nx5409, nx5411, 
         nx5413, nx5415, nx5417, nx5419, nx5421, nx5423, nx5425, nx5427, nx5429, 
         nx5431, nx5433, nx5435, nx5437, nx5439, nx5441, nx5443, nx5445, nx5447, 
         nx5449, nx5451, nx5453, nx5455, nx5457, nx5459, nx5461, nx5463, nx5465, 
         nx5467, nx5469, nx5471, nx5473, nx5475, nx5477, nx5479, nx5481, nx5483, 
         nx5485, nx5487, nx5489, nx5491, nx5493, nx5495, nx5501, nx5507, nx5511, 
         nx5517, nx5521, nx5525, nx5527, nx5531, nx5537, nx5539, nx5543, nx5547, 
         nx5549, nx5553, nx5559, nx5561, nx5563, nx5567, nx5569, nx5573, nx5581, 
         nx5585, nx5589, nx5591, nx5595, nx5601, nx5603, nx5607, nx5611, nx5613, 
         nx5617, nx5623, nx5625, nx5627, nx5631, nx5633, nx5637, nx5645, nx5649, 
         nx5653, nx5655, nx5659, nx5665, nx5667, nx5671, nx5675, nx5677, nx5681, 
         nx5687, nx5689, nx5691, nx5695, nx5697, nx5701, nx5709, nx5713, nx5717, 
         nx5719, nx5723, nx5729, nx5731, nx5735, nx5741, nx5745, nx5747, nx5749, 
         nx5755, nx5759, nx5763, nx5769, nx5773, nx5775, nx5777, nx5783, nx5787, 
         nx5791, nx5797, nx5801, nx5803, nx5805, nx5811, nx5815, nx5819, nx5825, 
         nx5829, nx5831, nx5833, nx5839, nx5843, nx5845, nx5849, nx5853, nx5855, 
         nx5857, nx5861, nx5863, nx5865, nx5867, nx5869, nx5871, nx5873, nx5877, 
         nx5879, nx5881, nx5883, nx5885, nx5887, nx5889, nx5893, nx5895, nx5897, 
         nx5899, nx5903, nx5905, nx5919, nx5929, nx5939, nx5949, nx5959, nx5963, 
         nx5967, nx5975, nx5981, nx5987, nx5989, nx5995, nx6001, nx6003, nx6011, 
         nx6013, nx6015, nx6017, nx6021, nx6033, nx6039, nx6041, nx6049, nx6051, 
         nx6053, nx6055, nx6059, nx6071, nx6077, nx6079, nx6087, nx6089, nx6091, 
         nx6093, nx6097, nx6109, nx6115, nx6117, nx6125, nx6127, nx6129, nx6131, 
         nx6135, nx6147, nx6153, nx6155, nx6163, nx6165, nx6167, nx6169, nx6173, 
         nx6185, nx6191, nx6193, nx6201, nx6203, nx6205, nx6207, nx6211, nx6223, 
         nx6229, nx6231, nx6239, nx6241, nx6243, nx6247, nx6251, nx6255, nx6257, 
         nx6261, nx6265, nx6267, nx6271, nx6279, nx6285, nx6293, nx6297, nx6303, 
         nx6307, nx6314, nx6316, nx6371, nx6373, nx6375, nx6377, nx6379, nx6381, 
         nx6383, nx6385, nx6387, nx6389, nx6391, nx6393, nx6395, nx6397, nx6399, 
         nx6401, nx6403, nx6405, nx6407, nx6409, nx6411, nx6413, nx6415, nx6417, 
         nx6419, nx6421, nx6423, nx6425, nx6427, nx6429, nx6431, nx6433, nx6435, 
         nx6437, nx6441, nx6447, nx6453, nx6460, nx6462, nx6464, nx6466, nx6468, 
         nx6470, nx6472, nx6475, nx6477, nx6479, nx6481, nx6483, nx6485, nx6487, 
         nx6489, nx6491;



    xnor2 ix1246 (.Y (nx1245), .A0 (nx1247), .A1 (nx1311)) ;
    xnor2 ix1248 (.Y (nx1247), .A0 (nx8694), .A1 (nx1303)) ;
    nor02ii ix8695 (.Y (nx8694), .A0 (nx1251), .A1 (nx8680)) ;
    xnor2 ix1252 (.Y (nx1251), .A0 (nx1253), .A1 (nx1281)) ;
    mux21_ni ix1254 (.Y (nx1253), .A0 (nx1255), .A1 (nx1277), .S0 (nx1279)) ;
    mux21_ni ix1256 (.Y (nx1255), .A0 (nx1257), .A1 (nx1273), .S0 (nx1275)) ;
    mux21_ni ix1258 (.Y (nx1257), .A0 (nx1259), .A1 (nx1269), .S0 (nx1271)) ;
    mux21_ni ix1260 (.Y (nx1259), .A0 (nx1261), .A1 (nx1265), .S0 (nx1267)) ;
    aoi32 ix1262 (.Y (nx1261), .A0 (input_b[23]), .A1 (input_a[23]), .A2 (nx8620
          ), .B0 (input_a[24]), .B1 (input_b[24])) ;
    inv02 ix1266 (.Y (nx1265), .A (input_a[25])) ;
    xnor2 ix1268 (.Y (nx1267), .A0 (input_b[25]), .A1 (input_a[25])) ;
    inv02 ix1270 (.Y (nx1269), .A (input_a[26])) ;
    xnor2 ix1272 (.Y (nx1271), .A0 (input_b[26]), .A1 (input_a[26])) ;
    inv02 ix1274 (.Y (nx1273), .A (input_a[27])) ;
    xnor2 ix1276 (.Y (nx1275), .A0 (input_b[27]), .A1 (input_a[27])) ;
    inv02 ix1278 (.Y (nx1277), .A (input_a[28])) ;
    xnor2 ix1280 (.Y (nx1279), .A0 (input_b[28]), .A1 (input_a[28])) ;
    xnor2 ix1282 (.Y (nx1281), .A0 (input_b[29]), .A1 (input_a[29])) ;
    nor02ii ix8681 (.Y (nx8680), .A0 (nx1285), .A1 (nx8666)) ;
    xnor2 ix1286 (.Y (nx1285), .A0 (nx1255), .A1 (nx1279)) ;
    nor02ii ix8667 (.Y (nx8666), .A0 (nx1289), .A1 (nx8652)) ;
    xnor2 ix1290 (.Y (nx1289), .A0 (nx1257), .A1 (nx1275)) ;
    nor02ii ix8653 (.Y (nx8652), .A0 (nx1293), .A1 (nx6427)) ;
    xnor2 ix1294 (.Y (nx1293), .A0 (nx1259), .A1 (nx1271)) ;
    nor04 ix8639 (.Y (nx8638), .A0 (nx8604), .A1 (nx1299), .A2 (nx1301), .A3 (
          nx1267)) ;
    nor02_2x ix1300 (.Y (nx1299), .A0 (input_a[23]), .A1 (input_b[23])) ;
    xnor2 ix1302 (.Y (nx1301), .A0 (input_b[24]), .A1 (input_a[24])) ;
    xnor2 ix1304 (.Y (nx1303), .A0 (nx1305), .A1 (nx1309)) ;
    mux21_ni ix1306 (.Y (nx1305), .A0 (nx1253), .A1 (nx1307), .S0 (nx1281)) ;
    inv02 ix1308 (.Y (nx1307), .A (input_a[29])) ;
    xnor2 ix1310 (.Y (nx1309), .A0 (input_a[30]), .A1 (input_b[30])) ;
    nand02_2x ix1312 (.Y (nx1311), .A0 (nx8714), .A1 (nx6431)) ;
    xnor2 ix8715 (.Y (nx8714), .A0 (nx8680), .A1 (nx1251)) ;
    nor02ii ix8755 (.Y (nx8754), .A0 (nx1317), .A1 (nx8720)) ;
    nand02_2x ix1318 (.Y (nx1317), .A0 (nx8726), .A1 (nx6429)) ;
    xnor2 ix8727 (.Y (nx8726), .A0 (nx8652), .A1 (nx1289)) ;
    nor02ii ix8751 (.Y (nx8750), .A0 (nx1323), .A1 (nx8732)) ;
    nand02_2x ix1324 (.Y (nx1323), .A0 (nx8738), .A1 (nx8746)) ;
    xnor2 ix8739 (.Y (nx8738), .A0 (nx8624), .A1 (nx1335)) ;
    nor02_2x ix8625 (.Y (nx8624), .A0 (nx1329), .A1 (nx1333)) ;
    oai21 ix1330 (.Y (nx1329), .A0 (input_a[23]), .A1 (input_b[23]), .B0 (nx1331
          )) ;
    nand02_2x ix1332 (.Y (nx1331), .A0 (input_b[23]), .A1 (input_a[23])) ;
    xnor2 ix1334 (.Y (nx1333), .A0 (nx1331), .A1 (nx1301)) ;
    xnor2 ix1336 (.Y (nx1335), .A0 (nx1261), .A1 (nx1267)) ;
    nor03_2x ix8747 (.Y (nx8746), .A0 (nx8610), .A1 (nx1333), .A2 (nx6491)) ;
    xnor2 ix1342 (.Y (nx1341), .A0 (nx1343), .A1 (nx5735)) ;
    nor02_2x ix1344 (.Y (nx1343), .A0 (nx7912), .A1 (nx4288)) ;
    mux21_ni ix7913 (.Y (nx7912), .A0 (nx4290), .A1 (nx7908), .S0 (nx4592)) ;
    aoi32 ix1350 (.Y (nx1349), .A0 (input_b[22]), .A1 (input_a[22]), .A2 (
          input_a[21]), .B0 (nx6389), .B1 (nx4030)) ;
    aoi32 ix1360 (.Y (nx1359), .A0 (input_b[22]), .A1 (input_a[20]), .A2 (
          input_a[19]), .B0 (nx6387), .B1 (nx4046)) ;
    aoi32 ix1368 (.Y (nx1367), .A0 (input_b[22]), .A1 (input_a[18]), .A2 (
          input_a[17]), .B0 (nx6385), .B1 (nx4062)) ;
    aoi32 ix1376 (.Y (nx1375), .A0 (input_b[22]), .A1 (input_a[16]), .A2 (
          input_a[15]), .B0 (nx6383), .B1 (nx4078)) ;
    aoi32 ix1384 (.Y (nx1383), .A0 (input_b[22]), .A1 (input_a[14]), .A2 (
          input_a[13]), .B0 (nx6381), .B1 (nx4094)) ;
    aoi32 ix1392 (.Y (nx1391), .A0 (input_b[22]), .A1 (input_a[12]), .A2 (
          input_a[11]), .B0 (nx6379), .B1 (nx4110)) ;
    aoi32 ix1400 (.Y (nx1399), .A0 (input_b[22]), .A1 (input_a[10]), .A2 (
          input_a[9]), .B0 (nx6377), .B1 (nx4126)) ;
    aoi32 ix1408 (.Y (nx1407), .A0 (input_b[22]), .A1 (input_a[8]), .A2 (
          input_a[7]), .B0 (nx6375), .B1 (nx4142)) ;
    aoi32 ix1416 (.Y (nx1415), .A0 (input_b[22]), .A1 (input_a[6]), .A2 (
          input_a[5]), .B0 (nx6373), .B1 (nx4158)) ;
    aoi32 ix1424 (.Y (nx1423), .A0 (input_b[22]), .A1 (input_a[4]), .A2 (
          input_a[3]), .B0 (nx6371), .B1 (nx4174)) ;
    ao21 ix1432 (.Y (nx1431), .A0 (nx1433), .A1 (nx1435), .B0 (nx6441)) ;
    nand02_2x ix1434 (.Y (nx1433), .A0 (input_b[22]), .A1 (input_a[0])) ;
    nand02_2x ix1436 (.Y (nx1435), .A0 (input_b[22]), .A1 (input_a[2])) ;
    nand02_2x ix1442 (.Y (nx1441), .A0 (input_b[22]), .A1 (input_a[3])) ;
    xnor2 ix4175 (.Y (nx4174), .A0 (input_a[3]), .A1 (nx1445)) ;
    nand02_2x ix1446 (.Y (nx1445), .A0 (input_b[22]), .A1 (input_a[4])) ;
    nand02_2x ix1450 (.Y (nx1449), .A0 (input_b[22]), .A1 (input_a[5])) ;
    xnor2 ix4159 (.Y (nx4158), .A0 (input_a[5]), .A1 (nx1453)) ;
    nand02_2x ix1454 (.Y (nx1453), .A0 (input_b[22]), .A1 (input_a[6])) ;
    nand02_2x ix1458 (.Y (nx1457), .A0 (input_b[22]), .A1 (input_a[7])) ;
    xnor2 ix4143 (.Y (nx4142), .A0 (input_a[7]), .A1 (nx1461)) ;
    nand02_2x ix1462 (.Y (nx1461), .A0 (input_b[22]), .A1 (input_a[8])) ;
    nand02_2x ix1466 (.Y (nx1465), .A0 (input_b[22]), .A1 (input_a[9])) ;
    xnor2 ix4127 (.Y (nx4126), .A0 (input_a[9]), .A1 (nx1469)) ;
    nand02_2x ix1470 (.Y (nx1469), .A0 (input_b[22]), .A1 (input_a[10])) ;
    nand02_2x ix1474 (.Y (nx1473), .A0 (input_b[22]), .A1 (input_a[11])) ;
    xnor2 ix4111 (.Y (nx4110), .A0 (input_a[11]), .A1 (nx1477)) ;
    nand02_2x ix1478 (.Y (nx1477), .A0 (input_b[22]), .A1 (input_a[12])) ;
    nand02_2x ix1482 (.Y (nx1481), .A0 (input_b[22]), .A1 (input_a[13])) ;
    xnor2 ix4095 (.Y (nx4094), .A0 (input_a[13]), .A1 (nx1485)) ;
    nand02_2x ix1486 (.Y (nx1485), .A0 (input_b[22]), .A1 (input_a[14])) ;
    nand02_2x ix1490 (.Y (nx1489), .A0 (input_b[22]), .A1 (input_a[15])) ;
    xnor2 ix4079 (.Y (nx4078), .A0 (input_a[15]), .A1 (nx1493)) ;
    nand02_2x ix1494 (.Y (nx1493), .A0 (input_b[22]), .A1 (input_a[16])) ;
    nand02_2x ix1498 (.Y (nx1497), .A0 (input_b[22]), .A1 (input_a[17])) ;
    xnor2 ix4063 (.Y (nx4062), .A0 (input_a[17]), .A1 (nx1501)) ;
    nand02_2x ix1502 (.Y (nx1501), .A0 (input_b[22]), .A1 (input_a[18])) ;
    nand02_2x ix1506 (.Y (nx1505), .A0 (input_b[22]), .A1 (input_a[19])) ;
    xnor2 ix4047 (.Y (nx4046), .A0 (input_a[19]), .A1 (nx1509)) ;
    nand02_2x ix1510 (.Y (nx1509), .A0 (input_b[22]), .A1 (input_a[20])) ;
    nand02_2x ix1514 (.Y (nx1513), .A0 (input_b[22]), .A1 (input_a[21])) ;
    xnor2 ix4031 (.Y (nx4030), .A0 (input_a[21]), .A1 (nx1517)) ;
    nand02_2x ix1518 (.Y (nx1517), .A0 (input_b[22]), .A1 (input_a[22])) ;
    oai21 ix1520 (.Y (nx1519), .A0 (input_a[22]), .A1 (input_b[22]), .B0 (nx1517
          )) ;
    mux21_ni ix7909 (.Y (nx7908), .A0 (nx7904), .A1 (nx4598), .S0 (nx5719)) ;
    xnor2 ix1526 (.Y (nx1525), .A0 (nx1527), .A1 (nx1889)) ;
    mux21_ni ix1528 (.Y (nx1527), .A0 (nx1529), .A1 (nx1875), .S0 (nx1877)) ;
    mux21_ni ix1530 (.Y (nx1529), .A0 (nx1531), .A1 (nx1533), .S0 (nx4622)) ;
    nand02_2x ix1532 (.Y (nx1531), .A0 (input_b[20]), .A1 (input_a[21])) ;
    mux21_ni ix1534 (.Y (nx1533), .A0 (nx1535), .A1 (nx1847), .S0 (nx1849)) ;
    mux21_ni ix1536 (.Y (nx1535), .A0 (nx1537), .A1 (nx1539), .S0 (nx4642)) ;
    nand02_2x ix1538 (.Y (nx1537), .A0 (input_b[20]), .A1 (input_a[19])) ;
    mux21_ni ix1540 (.Y (nx1539), .A0 (nx1541), .A1 (nx1819), .S0 (nx1821)) ;
    mux21_ni ix1542 (.Y (nx1541), .A0 (nx1543), .A1 (nx1545), .S0 (nx4662)) ;
    nand02_2x ix1544 (.Y (nx1543), .A0 (input_b[20]), .A1 (input_a[17])) ;
    mux21_ni ix1546 (.Y (nx1545), .A0 (nx1547), .A1 (nx1791), .S0 (nx1793)) ;
    mux21_ni ix1548 (.Y (nx1547), .A0 (nx1549), .A1 (nx1551), .S0 (nx4682)) ;
    nand02_2x ix1550 (.Y (nx1549), .A0 (input_b[20]), .A1 (input_a[15])) ;
    mux21_ni ix1552 (.Y (nx1551), .A0 (nx1553), .A1 (nx1763), .S0 (nx1765)) ;
    mux21_ni ix1554 (.Y (nx1553), .A0 (nx1555), .A1 (nx1557), .S0 (nx4702)) ;
    nand02_2x ix1556 (.Y (nx1555), .A0 (input_b[20]), .A1 (input_a[13])) ;
    mux21_ni ix1558 (.Y (nx1557), .A0 (nx1559), .A1 (nx1735), .S0 (nx1737)) ;
    mux21_ni ix1560 (.Y (nx1559), .A0 (nx1561), .A1 (nx1563), .S0 (nx4722)) ;
    nand02_2x ix1562 (.Y (nx1561), .A0 (input_b[20]), .A1 (input_a[11])) ;
    mux21_ni ix1564 (.Y (nx1563), .A0 (nx1565), .A1 (nx1707), .S0 (nx1709)) ;
    mux21_ni ix1566 (.Y (nx1565), .A0 (nx1567), .A1 (nx1569), .S0 (nx4742)) ;
    nand02_2x ix1568 (.Y (nx1567), .A0 (input_b[20]), .A1 (input_a[9])) ;
    mux21_ni ix1570 (.Y (nx1569), .A0 (nx1571), .A1 (nx1679), .S0 (nx1681)) ;
    mux21_ni ix1572 (.Y (nx1571), .A0 (nx1573), .A1 (nx1575), .S0 (nx4762)) ;
    nand02_2x ix1574 (.Y (nx1573), .A0 (input_b[20]), .A1 (input_a[7])) ;
    mux21_ni ix1576 (.Y (nx1575), .A0 (nx1577), .A1 (nx1651), .S0 (nx1653)) ;
    mux21_ni ix1578 (.Y (nx1577), .A0 (nx1579), .A1 (nx1581), .S0 (nx4782)) ;
    nand02_2x ix1580 (.Y (nx1579), .A0 (input_b[20]), .A1 (input_a[5])) ;
    mux21_ni ix1582 (.Y (nx1581), .A0 (nx1583), .A1 (nx1619), .S0 (nx1621)) ;
    mux21_ni ix1584 (.Y (nx1583), .A0 (nx1585), .A1 (nx1587), .S0 (nx3804)) ;
    nand02_2x ix1586 (.Y (nx1585), .A0 (input_b[20]), .A1 (input_a[3])) ;
    mux21_ni ix1588 (.Y (nx1587), .A0 (nx1589), .A1 (nx1591), .S0 (nx1593)) ;
    nand02_2x ix1592 (.Y (nx1591), .A0 (input_b[20]), .A1 (input_a[2])) ;
    xnor2 ix1594 (.Y (nx1593), .A0 (nx1595), .A1 (nx1591)) ;
    ao21 ix1596 (.Y (nx1595), .A0 (input_b[21]), .A1 (nx3190), .B0 (nx1601)) ;
    aoi22 ix1602 (.Y (nx1601), .A0 (input_b[22]), .A1 (input_a[0]), .B0 (
          input_b[21]), .B1 (input_a[1])) ;
    xnor2 ix3805 (.Y (nx3804), .A0 (nx3800), .A1 (nx1585)) ;
    xnor2 ix3801 (.Y (nx3800), .A0 (nx3192), .A1 (nx1611)) ;
    inv02 ix1610 (.Y (nx1609), .A (input_b[21])) ;
    xnor2 ix1612 (.Y (nx1611), .A0 (nx1613), .A1 (nx1617)) ;
    ao21 ix1614 (.Y (nx1613), .A0 (nx1615), .A1 (nx6447), .B0 (nx3190)) ;
    nand02_2x ix1616 (.Y (nx1615), .A0 (input_b[22]), .A1 (input_a[1])) ;
    nand02_2x ix1618 (.Y (nx1617), .A0 (input_b[21]), .A1 (input_a[2])) ;
    nand02_2x ix1620 (.Y (nx1619), .A0 (input_b[20]), .A1 (input_a[4])) ;
    xnor2 ix1622 (.Y (nx1621), .A0 (nx1623), .A1 (nx1619)) ;
    xnor2 ix1624 (.Y (nx1623), .A0 (nx1625), .A1 (nx1629)) ;
    aoi32 ix1626 (.Y (nx1625), .A0 (input_b[21]), .A1 (nx3190), .A2 (input_a[2])
          , .B0 (nx3796), .B1 (nx1611)) ;
    xnor2 ix1630 (.Y (nx1629), .A0 (nx1631), .A1 (nx1635)) ;
    xnor2 ix1632 (.Y (nx1631), .A0 (nx3190), .A1 (nx4190)) ;
    xnor2 ix4191 (.Y (nx4190), .A0 (input_a[1]), .A1 (nx1435)) ;
    nand02_2x ix1636 (.Y (nx1635), .A0 (input_b[21]), .A1 (input_a[3])) ;
    xnor2 ix4783 (.Y (nx4782), .A0 (nx4780), .A1 (nx1579)) ;
    xnor2 ix4781 (.Y (nx4780), .A0 (nx1641), .A1 (nx4484)) ;
    mux21_ni ix1642 (.Y (nx1641), .A0 (nx1625), .A1 (nx1635), .S0 (nx1629)) ;
    xnor2 ix4485 (.Y (nx4484), .A0 (nx4482), .A1 (nx1649)) ;
    xnor2 ix4483 (.Y (nx4482), .A0 (nx1431), .A1 (nx4182)) ;
    xnor2 ix4183 (.Y (nx4182), .A0 (input_a[2]), .A1 (nx1441)) ;
    nand02_2x ix1650 (.Y (nx1649), .A0 (input_b[21]), .A1 (input_a[4])) ;
    nand02_2x ix1652 (.Y (nx1651), .A0 (input_b[20]), .A1 (input_a[6])) ;
    xnor2 ix1654 (.Y (nx1653), .A0 (nx1655), .A1 (nx1651)) ;
    xnor2 ix1656 (.Y (nx1655), .A0 (nx1657), .A1 (nx1659)) ;
    mux21_ni ix1658 (.Y (nx1657), .A0 (nx1649), .A1 (nx1641), .S0 (nx4484)) ;
    xnor2 ix1660 (.Y (nx1659), .A0 (nx1661), .A1 (nx1663)) ;
    xnor2 ix1662 (.Y (nx1661), .A0 (nx6371), .A1 (nx4174)) ;
    nand02_2x ix1664 (.Y (nx1663), .A0 (input_b[21]), .A1 (input_a[5])) ;
    xnor2 ix4763 (.Y (nx4762), .A0 (nx4760), .A1 (nx1573)) ;
    xnor2 ix4761 (.Y (nx4760), .A0 (nx1669), .A1 (nx4464)) ;
    mux21_ni ix1670 (.Y (nx1669), .A0 (nx1657), .A1 (nx1663), .S0 (nx1659)) ;
    xnor2 ix4465 (.Y (nx4464), .A0 (nx4462), .A1 (nx1677)) ;
    xnor2 ix4463 (.Y (nx4462), .A0 (nx1423), .A1 (nx4166)) ;
    xnor2 ix4167 (.Y (nx4166), .A0 (input_a[4]), .A1 (nx1449)) ;
    nand02_2x ix1678 (.Y (nx1677), .A0 (input_b[21]), .A1 (input_a[6])) ;
    nand02_2x ix1680 (.Y (nx1679), .A0 (input_b[20]), .A1 (input_a[8])) ;
    xnor2 ix1682 (.Y (nx1681), .A0 (nx1683), .A1 (nx1679)) ;
    xnor2 ix1684 (.Y (nx1683), .A0 (nx1685), .A1 (nx1687)) ;
    mux21_ni ix1686 (.Y (nx1685), .A0 (nx1677), .A1 (nx1669), .S0 (nx4464)) ;
    xnor2 ix1688 (.Y (nx1687), .A0 (nx1689), .A1 (nx1691)) ;
    xnor2 ix1690 (.Y (nx1689), .A0 (nx6373), .A1 (nx4158)) ;
    nand02_2x ix1692 (.Y (nx1691), .A0 (input_b[21]), .A1 (input_a[7])) ;
    xnor2 ix4743 (.Y (nx4742), .A0 (nx4740), .A1 (nx1567)) ;
    xnor2 ix4741 (.Y (nx4740), .A0 (nx1697), .A1 (nx4444)) ;
    mux21_ni ix1698 (.Y (nx1697), .A0 (nx1685), .A1 (nx1691), .S0 (nx1687)) ;
    xnor2 ix4445 (.Y (nx4444), .A0 (nx4442), .A1 (nx1705)) ;
    xnor2 ix4443 (.Y (nx4442), .A0 (nx1415), .A1 (nx4150)) ;
    xnor2 ix4151 (.Y (nx4150), .A0 (input_a[6]), .A1 (nx1457)) ;
    nand02_2x ix1706 (.Y (nx1705), .A0 (input_b[21]), .A1 (input_a[8])) ;
    nand02_2x ix1708 (.Y (nx1707), .A0 (input_b[20]), .A1 (input_a[10])) ;
    xnor2 ix1710 (.Y (nx1709), .A0 (nx1711), .A1 (nx1707)) ;
    xnor2 ix1712 (.Y (nx1711), .A0 (nx1713), .A1 (nx1715)) ;
    mux21_ni ix1714 (.Y (nx1713), .A0 (nx1705), .A1 (nx1697), .S0 (nx4444)) ;
    xnor2 ix1716 (.Y (nx1715), .A0 (nx1717), .A1 (nx1719)) ;
    xnor2 ix1718 (.Y (nx1717), .A0 (nx6375), .A1 (nx4142)) ;
    nand02_2x ix1720 (.Y (nx1719), .A0 (input_b[21]), .A1 (input_a[9])) ;
    xnor2 ix4723 (.Y (nx4722), .A0 (nx4720), .A1 (nx1561)) ;
    xnor2 ix4721 (.Y (nx4720), .A0 (nx1725), .A1 (nx4424)) ;
    mux21_ni ix1726 (.Y (nx1725), .A0 (nx1713), .A1 (nx1719), .S0 (nx1715)) ;
    xnor2 ix4425 (.Y (nx4424), .A0 (nx4422), .A1 (nx1733)) ;
    xnor2 ix4423 (.Y (nx4422), .A0 (nx1407), .A1 (nx4134)) ;
    xnor2 ix4135 (.Y (nx4134), .A0 (input_a[8]), .A1 (nx1465)) ;
    nand02_2x ix1734 (.Y (nx1733), .A0 (input_b[21]), .A1 (input_a[10])) ;
    nand02_2x ix1736 (.Y (nx1735), .A0 (input_b[20]), .A1 (input_a[12])) ;
    xnor2 ix1738 (.Y (nx1737), .A0 (nx1739), .A1 (nx1735)) ;
    xnor2 ix1740 (.Y (nx1739), .A0 (nx1741), .A1 (nx1743)) ;
    mux21_ni ix1742 (.Y (nx1741), .A0 (nx1733), .A1 (nx1725), .S0 (nx4424)) ;
    xnor2 ix1744 (.Y (nx1743), .A0 (nx1745), .A1 (nx1747)) ;
    xnor2 ix1746 (.Y (nx1745), .A0 (nx6377), .A1 (nx4126)) ;
    nand02_2x ix1748 (.Y (nx1747), .A0 (input_b[21]), .A1 (input_a[11])) ;
    xnor2 ix4703 (.Y (nx4702), .A0 (nx4700), .A1 (nx1555)) ;
    xnor2 ix4701 (.Y (nx4700), .A0 (nx1753), .A1 (nx4404)) ;
    mux21_ni ix1754 (.Y (nx1753), .A0 (nx1741), .A1 (nx1747), .S0 (nx1743)) ;
    xnor2 ix4405 (.Y (nx4404), .A0 (nx4402), .A1 (nx1761)) ;
    xnor2 ix4403 (.Y (nx4402), .A0 (nx1399), .A1 (nx4118)) ;
    xnor2 ix4119 (.Y (nx4118), .A0 (input_a[10]), .A1 (nx1473)) ;
    nand02_2x ix1762 (.Y (nx1761), .A0 (input_b[21]), .A1 (input_a[12])) ;
    nand02_2x ix1764 (.Y (nx1763), .A0 (input_b[20]), .A1 (input_a[14])) ;
    xnor2 ix1766 (.Y (nx1765), .A0 (nx1767), .A1 (nx1763)) ;
    xnor2 ix1768 (.Y (nx1767), .A0 (nx1769), .A1 (nx1771)) ;
    mux21_ni ix1770 (.Y (nx1769), .A0 (nx1761), .A1 (nx1753), .S0 (nx4404)) ;
    xnor2 ix1772 (.Y (nx1771), .A0 (nx1773), .A1 (nx1775)) ;
    xnor2 ix1774 (.Y (nx1773), .A0 (nx6379), .A1 (nx4110)) ;
    nand02_2x ix1776 (.Y (nx1775), .A0 (input_b[21]), .A1 (input_a[13])) ;
    xnor2 ix4683 (.Y (nx4682), .A0 (nx4680), .A1 (nx1549)) ;
    xnor2 ix4681 (.Y (nx4680), .A0 (nx1781), .A1 (nx4384)) ;
    mux21_ni ix1782 (.Y (nx1781), .A0 (nx1769), .A1 (nx1775), .S0 (nx1771)) ;
    xnor2 ix4385 (.Y (nx4384), .A0 (nx4382), .A1 (nx1789)) ;
    xnor2 ix4383 (.Y (nx4382), .A0 (nx1391), .A1 (nx4102)) ;
    xnor2 ix4103 (.Y (nx4102), .A0 (input_a[12]), .A1 (nx1481)) ;
    nand02_2x ix1790 (.Y (nx1789), .A0 (input_b[21]), .A1 (input_a[14])) ;
    nand02_2x ix1792 (.Y (nx1791), .A0 (input_b[20]), .A1 (input_a[16])) ;
    xnor2 ix1794 (.Y (nx1793), .A0 (nx1795), .A1 (nx1791)) ;
    xnor2 ix1796 (.Y (nx1795), .A0 (nx1797), .A1 (nx1799)) ;
    mux21_ni ix1798 (.Y (nx1797), .A0 (nx1789), .A1 (nx1781), .S0 (nx4384)) ;
    xnor2 ix1800 (.Y (nx1799), .A0 (nx1801), .A1 (nx1803)) ;
    xnor2 ix1802 (.Y (nx1801), .A0 (nx6381), .A1 (nx4094)) ;
    nand02_2x ix1804 (.Y (nx1803), .A0 (input_b[21]), .A1 (input_a[15])) ;
    xnor2 ix4663 (.Y (nx4662), .A0 (nx4660), .A1 (nx1543)) ;
    xnor2 ix4661 (.Y (nx4660), .A0 (nx1809), .A1 (nx4364)) ;
    mux21_ni ix1810 (.Y (nx1809), .A0 (nx1797), .A1 (nx1803), .S0 (nx1799)) ;
    xnor2 ix4365 (.Y (nx4364), .A0 (nx4362), .A1 (nx1817)) ;
    xnor2 ix4363 (.Y (nx4362), .A0 (nx1383), .A1 (nx4086)) ;
    xnor2 ix4087 (.Y (nx4086), .A0 (input_a[14]), .A1 (nx1489)) ;
    nand02_2x ix1818 (.Y (nx1817), .A0 (input_b[21]), .A1 (input_a[16])) ;
    nand02_2x ix1820 (.Y (nx1819), .A0 (input_b[20]), .A1 (input_a[18])) ;
    xnor2 ix1822 (.Y (nx1821), .A0 (nx1823), .A1 (nx1819)) ;
    xnor2 ix1824 (.Y (nx1823), .A0 (nx1825), .A1 (nx1827)) ;
    mux21_ni ix1826 (.Y (nx1825), .A0 (nx1817), .A1 (nx1809), .S0 (nx4364)) ;
    xnor2 ix1828 (.Y (nx1827), .A0 (nx1829), .A1 (nx1831)) ;
    xnor2 ix1830 (.Y (nx1829), .A0 (nx6383), .A1 (nx4078)) ;
    nand02_2x ix1832 (.Y (nx1831), .A0 (input_b[21]), .A1 (input_a[17])) ;
    xnor2 ix4643 (.Y (nx4642), .A0 (nx4640), .A1 (nx1537)) ;
    xnor2 ix4641 (.Y (nx4640), .A0 (nx1837), .A1 (nx4344)) ;
    mux21_ni ix1838 (.Y (nx1837), .A0 (nx1825), .A1 (nx1831), .S0 (nx1827)) ;
    xnor2 ix4345 (.Y (nx4344), .A0 (nx4342), .A1 (nx1845)) ;
    xnor2 ix4343 (.Y (nx4342), .A0 (nx1375), .A1 (nx4070)) ;
    xnor2 ix4071 (.Y (nx4070), .A0 (input_a[16]), .A1 (nx1497)) ;
    nand02_2x ix1846 (.Y (nx1845), .A0 (input_b[21]), .A1 (input_a[18])) ;
    nand02_2x ix1848 (.Y (nx1847), .A0 (input_b[20]), .A1 (input_a[20])) ;
    xnor2 ix1850 (.Y (nx1849), .A0 (nx1851), .A1 (nx1847)) ;
    xnor2 ix1852 (.Y (nx1851), .A0 (nx1853), .A1 (nx1855)) ;
    mux21_ni ix1854 (.Y (nx1853), .A0 (nx1845), .A1 (nx1837), .S0 (nx4344)) ;
    xnor2 ix1856 (.Y (nx1855), .A0 (nx1857), .A1 (nx1859)) ;
    xnor2 ix1858 (.Y (nx1857), .A0 (nx6385), .A1 (nx4062)) ;
    nand02_2x ix1860 (.Y (nx1859), .A0 (input_b[21]), .A1 (input_a[19])) ;
    xnor2 ix4623 (.Y (nx4622), .A0 (nx4620), .A1 (nx1531)) ;
    xnor2 ix4621 (.Y (nx4620), .A0 (nx1865), .A1 (nx4324)) ;
    mux21_ni ix1866 (.Y (nx1865), .A0 (nx1853), .A1 (nx1859), .S0 (nx1855)) ;
    xnor2 ix4325 (.Y (nx4324), .A0 (nx4322), .A1 (nx1873)) ;
    xnor2 ix4323 (.Y (nx4322), .A0 (nx1367), .A1 (nx4054)) ;
    xnor2 ix4055 (.Y (nx4054), .A0 (input_a[18]), .A1 (nx1505)) ;
    nand02_2x ix1874 (.Y (nx1873), .A0 (input_b[21]), .A1 (input_a[20])) ;
    nand02_2x ix1876 (.Y (nx1875), .A0 (input_b[20]), .A1 (input_a[22])) ;
    xnor2 ix1878 (.Y (nx1877), .A0 (nx1879), .A1 (nx1875)) ;
    xnor2 ix1880 (.Y (nx1879), .A0 (nx1881), .A1 (nx1883)) ;
    mux21_ni ix1882 (.Y (nx1881), .A0 (nx1873), .A1 (nx1865), .S0 (nx4324)) ;
    xnor2 ix1884 (.Y (nx1883), .A0 (nx1885), .A1 (nx1887)) ;
    xnor2 ix1886 (.Y (nx1885), .A0 (nx6387), .A1 (nx4046)) ;
    nand02_2x ix1888 (.Y (nx1887), .A0 (input_b[21]), .A1 (input_a[21])) ;
    xnor2 ix1890 (.Y (nx1889), .A0 (input_b[20]), .A1 (nx4600)) ;
    xnor2 ix4601 (.Y (nx4600), .A0 (nx1893), .A1 (nx4304)) ;
    mux21_ni ix1894 (.Y (nx1893), .A0 (nx1881), .A1 (nx1887), .S0 (nx1883)) ;
    xnor2 ix4305 (.Y (nx4304), .A0 (nx4302), .A1 (nx1901)) ;
    xnor2 ix4303 (.Y (nx4302), .A0 (nx1359), .A1 (nx4038)) ;
    xnor2 ix4039 (.Y (nx4038), .A0 (input_a[20]), .A1 (nx1513)) ;
    nand02_2x ix1902 (.Y (nx1901), .A0 (input_b[21]), .A1 (input_a[22])) ;
    mux21_ni ix1904 (.Y (nx1903), .A0 (nx1905), .A1 (nx5689), .S0 (nx5697)) ;
    mux21_ni ix1906 (.Y (nx1905), .A0 (nx1907), .A1 (nx2263), .S0 (nx5684)) ;
    xnor2 ix1908 (.Y (nx1907), .A0 (nx1909), .A1 (nx2251)) ;
    mux21_ni ix1910 (.Y (nx1909), .A0 (nx1911), .A1 (nx2237), .S0 (nx2239)) ;
    mux21_ni ix1912 (.Y (nx1911), .A0 (nx1913), .A1 (nx1915), .S0 (nx5196)) ;
    nand02_2x ix1914 (.Y (nx1913), .A0 (input_b[18]), .A1 (input_a[21])) ;
    mux21_ni ix1916 (.Y (nx1915), .A0 (nx1917), .A1 (nx2211), .S0 (nx2213)) ;
    mux21_ni ix1918 (.Y (nx1917), .A0 (nx1919), .A1 (nx1921), .S0 (nx5216)) ;
    nand02_2x ix1920 (.Y (nx1919), .A0 (input_b[18]), .A1 (input_a[19])) ;
    mux21_ni ix1922 (.Y (nx1921), .A0 (nx1923), .A1 (nx2185), .S0 (nx2187)) ;
    mux21_ni ix1924 (.Y (nx1923), .A0 (nx1925), .A1 (nx1927), .S0 (nx5236)) ;
    nand02_2x ix1926 (.Y (nx1925), .A0 (input_b[18]), .A1 (input_a[17])) ;
    mux21_ni ix1928 (.Y (nx1927), .A0 (nx1929), .A1 (nx2159), .S0 (nx2161)) ;
    mux21_ni ix1930 (.Y (nx1929), .A0 (nx1931), .A1 (nx1933), .S0 (nx5256)) ;
    nand02_2x ix1932 (.Y (nx1931), .A0 (input_b[18]), .A1 (input_a[15])) ;
    mux21_ni ix1934 (.Y (nx1933), .A0 (nx1935), .A1 (nx2133), .S0 (nx2135)) ;
    mux21_ni ix1936 (.Y (nx1935), .A0 (nx1937), .A1 (nx1939), .S0 (nx5276)) ;
    nand02_2x ix1938 (.Y (nx1937), .A0 (input_b[18]), .A1 (input_a[13])) ;
    mux21_ni ix1940 (.Y (nx1939), .A0 (nx1941), .A1 (nx2107), .S0 (nx2109)) ;
    mux21_ni ix1942 (.Y (nx1941), .A0 (nx1943), .A1 (nx1945), .S0 (nx5296)) ;
    nand02_2x ix1944 (.Y (nx1943), .A0 (input_b[18]), .A1 (input_a[11])) ;
    mux21_ni ix1946 (.Y (nx1945), .A0 (nx1947), .A1 (nx2081), .S0 (nx2083)) ;
    mux21_ni ix1948 (.Y (nx1947), .A0 (nx1949), .A1 (nx1951), .S0 (nx5316)) ;
    nand02_2x ix1950 (.Y (nx1949), .A0 (input_b[18]), .A1 (input_a[9])) ;
    mux21_ni ix1952 (.Y (nx1951), .A0 (nx1953), .A1 (nx2055), .S0 (nx2057)) ;
    mux21_ni ix1954 (.Y (nx1953), .A0 (nx1955), .A1 (nx1957), .S0 (nx5336)) ;
    nand02_2x ix1956 (.Y (nx1955), .A0 (input_b[18]), .A1 (input_a[7])) ;
    mux21_ni ix1958 (.Y (nx1957), .A0 (nx1959), .A1 (nx2029), .S0 (nx2031)) ;
    mux21_ni ix1960 (.Y (nx1959), .A0 (nx1961), .A1 (nx1963), .S0 (nx3816)) ;
    nand02_2x ix1962 (.Y (nx1961), .A0 (input_b[18]), .A1 (input_a[5])) ;
    mux21_ni ix1964 (.Y (nx1963), .A0 (nx1965), .A1 (nx1967), .S0 (nx3218)) ;
    nand02_2x ix1966 (.Y (nx1965), .A0 (input_b[18]), .A1 (input_a[4])) ;
    mux21_ni ix1968 (.Y (nx1967), .A0 (nx1969), .A1 (nx1987), .S0 (nx1989)) ;
    mux21_ni ix1970 (.Y (nx1969), .A0 (nx1971), .A1 (nx1973), .S0 (nx2174)) ;
    nand02_2x ix1972 (.Y (nx1971), .A0 (input_b[18]), .A1 (input_a[2])) ;
    xnor2 ix2175 (.Y (nx2174), .A0 (nx2170), .A1 (nx1971)) ;
    inv02 ix1982 (.Y (nx1981), .A (input_b[19])) ;
    inv02 ix1984 (.Y (nx1983), .A (input_b[20])) ;
    aoi22 ix1986 (.Y (nx1985), .A0 (input_b[20]), .A1 (input_a[0]), .B0 (
          input_b[19]), .B1 (input_a[1])) ;
    nand02_2x ix1988 (.Y (nx1987), .A0 (input_b[18]), .A1 (input_a[3])) ;
    xnor2 ix1990 (.Y (nx1989), .A0 (nx1991), .A1 (nx1987)) ;
    xnor2 ix2663 (.Y (nx2662), .A0 (nx2658), .A1 (nx2001)) ;
    aoi22 ix2000 (.Y (nx1999), .A0 (input_b[21]), .A1 (input_a[0]), .B0 (
          input_b[20]), .B1 (input_a[1])) ;
    nand02_2x ix2002 (.Y (nx2001), .A0 (input_b[19]), .A1 (input_a[2])) ;
    xnor2 ix3219 (.Y (nx3218), .A0 (nx3214), .A1 (nx1965)) ;
    xnor2 ix3215 (.Y (nx3214), .A0 (nx2007), .A1 (nx3212)) ;
    mux21_ni ix2008 (.Y (nx2007), .A0 (nx2001), .A1 (nx2009), .S0 (nx2662)) ;
    xnor2 ix3213 (.Y (nx3212), .A0 (nx3208), .A1 (nx2015)) ;
    nand02_2x ix2016 (.Y (nx2015), .A0 (input_b[19]), .A1 (input_a[3])) ;
    xnor2 ix3817 (.Y (nx3816), .A0 (nx3812), .A1 (nx1961)) ;
    xnor2 ix3813 (.Y (nx3812), .A0 (nx2021), .A1 (nx3810)) ;
    mux21_ni ix2022 (.Y (nx2021), .A0 (nx2015), .A1 (nx2007), .S0 (nx3212)) ;
    xnor2 ix3811 (.Y (nx3810), .A0 (nx3806), .A1 (nx2027)) ;
    xnor2 ix3807 (.Y (nx3806), .A0 (nx1587), .A1 (nx3804)) ;
    nand02_2x ix2028 (.Y (nx2027), .A0 (input_b[19]), .A1 (input_a[4])) ;
    nand02_2x ix2030 (.Y (nx2029), .A0 (input_b[18]), .A1 (input_a[6])) ;
    xnor2 ix2032 (.Y (nx2031), .A0 (nx2033), .A1 (nx2029)) ;
    xnor2 ix2034 (.Y (nx2033), .A0 (nx2035), .A1 (nx2037)) ;
    mux21_ni ix2036 (.Y (nx2035), .A0 (nx2027), .A1 (nx2021), .S0 (nx3810)) ;
    xnor2 ix2038 (.Y (nx2037), .A0 (nx2039), .A1 (nx2041)) ;
    xnor2 ix2040 (.Y (nx2039), .A0 (nx1583), .A1 (nx1621)) ;
    nand02_2x ix2042 (.Y (nx2041), .A0 (input_b[19]), .A1 (input_a[5])) ;
    xnor2 ix5337 (.Y (nx5336), .A0 (nx5334), .A1 (nx1955)) ;
    xnor2 ix5335 (.Y (nx5334), .A0 (nx2047), .A1 (nx5066)) ;
    mux21_ni ix2048 (.Y (nx2047), .A0 (nx2035), .A1 (nx2041), .S0 (nx2037)) ;
    xnor2 ix5067 (.Y (nx5066), .A0 (nx5064), .A1 (nx2053)) ;
    xnor2 ix5065 (.Y (nx5064), .A0 (nx1581), .A1 (nx4782)) ;
    nand02_2x ix2054 (.Y (nx2053), .A0 (input_b[19]), .A1 (input_a[6])) ;
    nand02_2x ix2056 (.Y (nx2055), .A0 (input_b[18]), .A1 (input_a[8])) ;
    xnor2 ix2058 (.Y (nx2057), .A0 (nx2059), .A1 (nx2055)) ;
    xnor2 ix2060 (.Y (nx2059), .A0 (nx2061), .A1 (nx2063)) ;
    mux21_ni ix2062 (.Y (nx2061), .A0 (nx2053), .A1 (nx2047), .S0 (nx5066)) ;
    xnor2 ix2064 (.Y (nx2063), .A0 (nx2065), .A1 (nx2067)) ;
    xnor2 ix2066 (.Y (nx2065), .A0 (nx1577), .A1 (nx1653)) ;
    nand02_2x ix2068 (.Y (nx2067), .A0 (input_b[19]), .A1 (input_a[7])) ;
    xnor2 ix5317 (.Y (nx5316), .A0 (nx5314), .A1 (nx1949)) ;
    xnor2 ix5315 (.Y (nx5314), .A0 (nx2073), .A1 (nx5046)) ;
    mux21_ni ix2074 (.Y (nx2073), .A0 (nx2061), .A1 (nx2067), .S0 (nx2063)) ;
    xnor2 ix5047 (.Y (nx5046), .A0 (nx5044), .A1 (nx2079)) ;
    xnor2 ix5045 (.Y (nx5044), .A0 (nx1575), .A1 (nx4762)) ;
    nand02_2x ix2080 (.Y (nx2079), .A0 (input_b[19]), .A1 (input_a[8])) ;
    nand02_2x ix2082 (.Y (nx2081), .A0 (input_b[18]), .A1 (input_a[10])) ;
    xnor2 ix2084 (.Y (nx2083), .A0 (nx2085), .A1 (nx2081)) ;
    xnor2 ix2086 (.Y (nx2085), .A0 (nx2087), .A1 (nx2089)) ;
    mux21_ni ix2088 (.Y (nx2087), .A0 (nx2079), .A1 (nx2073), .S0 (nx5046)) ;
    xnor2 ix2090 (.Y (nx2089), .A0 (nx2091), .A1 (nx2093)) ;
    xnor2 ix2092 (.Y (nx2091), .A0 (nx1571), .A1 (nx1681)) ;
    nand02_2x ix2094 (.Y (nx2093), .A0 (input_b[19]), .A1 (input_a[9])) ;
    xnor2 ix5297 (.Y (nx5296), .A0 (nx5294), .A1 (nx1943)) ;
    xnor2 ix5295 (.Y (nx5294), .A0 (nx2099), .A1 (nx5026)) ;
    mux21_ni ix2100 (.Y (nx2099), .A0 (nx2087), .A1 (nx2093), .S0 (nx2089)) ;
    xnor2 ix5027 (.Y (nx5026), .A0 (nx5024), .A1 (nx2105)) ;
    xnor2 ix5025 (.Y (nx5024), .A0 (nx1569), .A1 (nx4742)) ;
    nand02_2x ix2106 (.Y (nx2105), .A0 (input_b[19]), .A1 (input_a[10])) ;
    nand02_2x ix2108 (.Y (nx2107), .A0 (input_b[18]), .A1 (input_a[12])) ;
    xnor2 ix2110 (.Y (nx2109), .A0 (nx2111), .A1 (nx2107)) ;
    xnor2 ix2112 (.Y (nx2111), .A0 (nx2113), .A1 (nx2115)) ;
    mux21_ni ix2114 (.Y (nx2113), .A0 (nx2105), .A1 (nx2099), .S0 (nx5026)) ;
    xnor2 ix2116 (.Y (nx2115), .A0 (nx2117), .A1 (nx2119)) ;
    xnor2 ix2118 (.Y (nx2117), .A0 (nx1565), .A1 (nx1709)) ;
    nand02_2x ix2120 (.Y (nx2119), .A0 (input_b[19]), .A1 (input_a[11])) ;
    xnor2 ix5277 (.Y (nx5276), .A0 (nx5274), .A1 (nx1937)) ;
    xnor2 ix5275 (.Y (nx5274), .A0 (nx2125), .A1 (nx5006)) ;
    mux21_ni ix2126 (.Y (nx2125), .A0 (nx2113), .A1 (nx2119), .S0 (nx2115)) ;
    xnor2 ix5007 (.Y (nx5006), .A0 (nx5004), .A1 (nx2131)) ;
    xnor2 ix5005 (.Y (nx5004), .A0 (nx1563), .A1 (nx4722)) ;
    nand02_2x ix2132 (.Y (nx2131), .A0 (input_b[19]), .A1 (input_a[12])) ;
    nand02_2x ix2134 (.Y (nx2133), .A0 (input_b[18]), .A1 (input_a[14])) ;
    xnor2 ix2136 (.Y (nx2135), .A0 (nx2137), .A1 (nx2133)) ;
    xnor2 ix2138 (.Y (nx2137), .A0 (nx2139), .A1 (nx2141)) ;
    mux21_ni ix2140 (.Y (nx2139), .A0 (nx2131), .A1 (nx2125), .S0 (nx5006)) ;
    xnor2 ix2142 (.Y (nx2141), .A0 (nx2143), .A1 (nx2145)) ;
    xnor2 ix2144 (.Y (nx2143), .A0 (nx1559), .A1 (nx1737)) ;
    nand02_2x ix2146 (.Y (nx2145), .A0 (input_b[19]), .A1 (input_a[13])) ;
    xnor2 ix5257 (.Y (nx5256), .A0 (nx5254), .A1 (nx1931)) ;
    xnor2 ix5255 (.Y (nx5254), .A0 (nx2151), .A1 (nx4986)) ;
    mux21_ni ix2152 (.Y (nx2151), .A0 (nx2139), .A1 (nx2145), .S0 (nx2141)) ;
    xnor2 ix4987 (.Y (nx4986), .A0 (nx4984), .A1 (nx2157)) ;
    xnor2 ix4985 (.Y (nx4984), .A0 (nx1557), .A1 (nx4702)) ;
    nand02_2x ix2158 (.Y (nx2157), .A0 (input_b[19]), .A1 (input_a[14])) ;
    nand02_2x ix2160 (.Y (nx2159), .A0 (input_b[18]), .A1 (input_a[16])) ;
    xnor2 ix2162 (.Y (nx2161), .A0 (nx2163), .A1 (nx2159)) ;
    xnor2 ix2164 (.Y (nx2163), .A0 (nx2165), .A1 (nx2167)) ;
    mux21_ni ix2166 (.Y (nx2165), .A0 (nx2157), .A1 (nx2151), .S0 (nx4986)) ;
    xnor2 ix2168 (.Y (nx2167), .A0 (nx2169), .A1 (nx2171)) ;
    xnor2 ix2170 (.Y (nx2169), .A0 (nx1553), .A1 (nx1765)) ;
    nand02_2x ix2172 (.Y (nx2171), .A0 (input_b[19]), .A1 (input_a[15])) ;
    xnor2 ix5237 (.Y (nx5236), .A0 (nx5234), .A1 (nx1925)) ;
    xnor2 ix5235 (.Y (nx5234), .A0 (nx2177), .A1 (nx4966)) ;
    mux21_ni ix2178 (.Y (nx2177), .A0 (nx2165), .A1 (nx2171), .S0 (nx2167)) ;
    xnor2 ix4967 (.Y (nx4966), .A0 (nx4964), .A1 (nx2183)) ;
    xnor2 ix4965 (.Y (nx4964), .A0 (nx1551), .A1 (nx4682)) ;
    nand02_2x ix2184 (.Y (nx2183), .A0 (input_b[19]), .A1 (input_a[16])) ;
    nand02_2x ix2186 (.Y (nx2185), .A0 (input_b[18]), .A1 (input_a[18])) ;
    xnor2 ix2188 (.Y (nx2187), .A0 (nx2189), .A1 (nx2185)) ;
    xnor2 ix2190 (.Y (nx2189), .A0 (nx2191), .A1 (nx2193)) ;
    mux21_ni ix2192 (.Y (nx2191), .A0 (nx2183), .A1 (nx2177), .S0 (nx4966)) ;
    xnor2 ix2194 (.Y (nx2193), .A0 (nx2195), .A1 (nx2197)) ;
    xnor2 ix2196 (.Y (nx2195), .A0 (nx1547), .A1 (nx1793)) ;
    nand02_2x ix2198 (.Y (nx2197), .A0 (input_b[19]), .A1 (input_a[17])) ;
    xnor2 ix5217 (.Y (nx5216), .A0 (nx5214), .A1 (nx1919)) ;
    xnor2 ix5215 (.Y (nx5214), .A0 (nx2203), .A1 (nx4946)) ;
    mux21_ni ix2204 (.Y (nx2203), .A0 (nx2191), .A1 (nx2197), .S0 (nx2193)) ;
    xnor2 ix4947 (.Y (nx4946), .A0 (nx4944), .A1 (nx2209)) ;
    xnor2 ix4945 (.Y (nx4944), .A0 (nx1545), .A1 (nx4662)) ;
    nand02_2x ix2210 (.Y (nx2209), .A0 (input_b[19]), .A1 (input_a[18])) ;
    nand02_2x ix2212 (.Y (nx2211), .A0 (input_b[18]), .A1 (input_a[20])) ;
    xnor2 ix2214 (.Y (nx2213), .A0 (nx2215), .A1 (nx2211)) ;
    xnor2 ix2216 (.Y (nx2215), .A0 (nx2217), .A1 (nx2219)) ;
    mux21_ni ix2218 (.Y (nx2217), .A0 (nx2209), .A1 (nx2203), .S0 (nx4946)) ;
    xnor2 ix2220 (.Y (nx2219), .A0 (nx2221), .A1 (nx2223)) ;
    xnor2 ix2222 (.Y (nx2221), .A0 (nx1541), .A1 (nx1821)) ;
    nand02_2x ix2224 (.Y (nx2223), .A0 (input_b[19]), .A1 (input_a[19])) ;
    xnor2 ix5197 (.Y (nx5196), .A0 (nx5194), .A1 (nx1913)) ;
    xnor2 ix5195 (.Y (nx5194), .A0 (nx2229), .A1 (nx4926)) ;
    mux21_ni ix2230 (.Y (nx2229), .A0 (nx2217), .A1 (nx2223), .S0 (nx2219)) ;
    xnor2 ix4927 (.Y (nx4926), .A0 (nx4924), .A1 (nx2235)) ;
    xnor2 ix4925 (.Y (nx4924), .A0 (nx1539), .A1 (nx4642)) ;
    nand02_2x ix2236 (.Y (nx2235), .A0 (input_b[19]), .A1 (input_a[20])) ;
    nand02_2x ix2238 (.Y (nx2237), .A0 (input_b[18]), .A1 (input_a[22])) ;
    xnor2 ix2240 (.Y (nx2239), .A0 (nx2241), .A1 (nx2237)) ;
    xnor2 ix2242 (.Y (nx2241), .A0 (nx2243), .A1 (nx2245)) ;
    mux21_ni ix2244 (.Y (nx2243), .A0 (nx2235), .A1 (nx2229), .S0 (nx4926)) ;
    xnor2 ix2246 (.Y (nx2245), .A0 (nx2247), .A1 (nx2249)) ;
    xnor2 ix2248 (.Y (nx2247), .A0 (nx1535), .A1 (nx1849)) ;
    nand02_2x ix2250 (.Y (nx2249), .A0 (input_b[19]), .A1 (input_a[21])) ;
    xnor2 ix2252 (.Y (nx2251), .A0 (input_b[18]), .A1 (nx5174)) ;
    xnor2 ix5175 (.Y (nx5174), .A0 (nx2255), .A1 (nx4906)) ;
    mux21_ni ix2256 (.Y (nx2255), .A0 (nx2243), .A1 (nx2249), .S0 (nx2245)) ;
    xnor2 ix4907 (.Y (nx4906), .A0 (nx4904), .A1 (nx2261)) ;
    xnor2 ix4905 (.Y (nx4904), .A0 (nx1533), .A1 (nx4622)) ;
    nand02_2x ix2262 (.Y (nx2261), .A0 (input_b[19]), .A1 (input_a[22])) ;
    mux21_ni ix7889 (.Y (nx7888), .A0 (nx5928), .A1 (nx7884), .S0 (nx6146)) ;
    mux21_ni ix2270 (.Y (nx2269), .A0 (nx2271), .A1 (nx2597), .S0 (nx2599)) ;
    mux21_ni ix2272 (.Y (nx2271), .A0 (nx2273), .A1 (nx2275), .S0 (nx5714)) ;
    nand02_2x ix2274 (.Y (nx2273), .A0 (input_b[16]), .A1 (input_a[21])) ;
    mux21_ni ix2276 (.Y (nx2275), .A0 (nx2277), .A1 (nx2571), .S0 (nx2573)) ;
    mux21_ni ix2278 (.Y (nx2277), .A0 (nx2279), .A1 (nx2281), .S0 (nx5734)) ;
    nand02_2x ix2280 (.Y (nx2279), .A0 (input_b[16]), .A1 (input_a[19])) ;
    mux21_ni ix2282 (.Y (nx2281), .A0 (nx2283), .A1 (nx2545), .S0 (nx2547)) ;
    mux21_ni ix2284 (.Y (nx2283), .A0 (nx2285), .A1 (nx2287), .S0 (nx5754)) ;
    nand02_2x ix2286 (.Y (nx2285), .A0 (input_b[16]), .A1 (input_a[17])) ;
    mux21_ni ix2288 (.Y (nx2287), .A0 (nx2289), .A1 (nx2519), .S0 (nx2521)) ;
    mux21_ni ix2290 (.Y (nx2289), .A0 (nx2291), .A1 (nx2293), .S0 (nx5774)) ;
    nand02_2x ix2292 (.Y (nx2291), .A0 (input_b[16]), .A1 (input_a[15])) ;
    mux21_ni ix2294 (.Y (nx2293), .A0 (nx2295), .A1 (nx2493), .S0 (nx2495)) ;
    mux21_ni ix2296 (.Y (nx2295), .A0 (nx2297), .A1 (nx2299), .S0 (nx5794)) ;
    nand02_2x ix2298 (.Y (nx2297), .A0 (input_b[16]), .A1 (input_a[13])) ;
    mux21_ni ix2300 (.Y (nx2299), .A0 (nx2301), .A1 (nx2467), .S0 (nx2469)) ;
    mux21_ni ix2302 (.Y (nx2301), .A0 (nx2303), .A1 (nx2305), .S0 (nx5814)) ;
    nand02_2x ix2304 (.Y (nx2303), .A0 (input_b[16]), .A1 (input_a[11])) ;
    mux21_ni ix2306 (.Y (nx2305), .A0 (nx2307), .A1 (nx2441), .S0 (nx2443)) ;
    mux21_ni ix2308 (.Y (nx2307), .A0 (nx2309), .A1 (nx2311), .S0 (nx5834)) ;
    nand02_2x ix2310 (.Y (nx2309), .A0 (input_b[16]), .A1 (input_a[9])) ;
    mux21_ni ix2312 (.Y (nx2311), .A0 (nx2313), .A1 (nx2415), .S0 (nx2417)) ;
    mux21_ni ix2314 (.Y (nx2313), .A0 (nx2315), .A1 (nx2317), .S0 (nx3828)) ;
    nand02_2x ix2316 (.Y (nx2315), .A0 (input_b[16]), .A1 (input_a[7])) ;
    mux21_ni ix2318 (.Y (nx2317), .A0 (nx2319), .A1 (nx2321), .S0 (nx3230)) ;
    nand02_2x ix2320 (.Y (nx2319), .A0 (input_b[16]), .A1 (input_a[6])) ;
    mux21_ni ix2322 (.Y (nx2321), .A0 (nx2323), .A1 (nx2377), .S0 (nx2379)) ;
    mux21_ni ix2324 (.Y (nx2323), .A0 (nx2325), .A1 (nx2361), .S0 (nx2363)) ;
    mux21_ni ix2326 (.Y (nx2325), .A0 (nx2327), .A1 (nx2345), .S0 (nx2347)) ;
    mux21_ni ix2328 (.Y (nx2327), .A0 (nx2329), .A1 (nx2331), .S0 (nx1366)) ;
    nand02_2x ix2330 (.Y (nx2329), .A0 (input_b[16]), .A1 (input_a[2])) ;
    xnor2 ix1367 (.Y (nx1366), .A0 (nx1362), .A1 (nx2329)) ;
    inv02 ix2340 (.Y (nx2339), .A (input_b[17])) ;
    inv02 ix2342 (.Y (nx2341), .A (input_b[18])) ;
    aoi22 ix2344 (.Y (nx2343), .A0 (input_b[18]), .A1 (input_a[0]), .B0 (
          input_b[17]), .B1 (input_a[1])) ;
    nand02_2x ix2346 (.Y (nx2345), .A0 (input_b[16]), .A1 (input_a[3])) ;
    xnor2 ix2348 (.Y (nx2347), .A0 (nx2349), .A1 (nx2345)) ;
    xnor2 ix1743 (.Y (nx1742), .A0 (nx1738), .A1 (nx2359)) ;
    aoi22 ix2358 (.Y (nx2357), .A0 (input_b[19]), .A1 (input_a[0]), .B0 (
          input_b[18]), .B1 (input_a[1])) ;
    nand02_2x ix2360 (.Y (nx2359), .A0 (input_b[17]), .A1 (input_a[2])) ;
    nand02_2x ix2362 (.Y (nx2361), .A0 (input_b[16]), .A1 (input_a[4])) ;
    xnor2 ix2364 (.Y (nx2363), .A0 (nx2365), .A1 (nx2361)) ;
    xnor2 ix2366 (.Y (nx2365), .A0 (nx2367), .A1 (nx2371)) ;
    mux21_ni ix2368 (.Y (nx2367), .A0 (nx2359), .A1 (nx2369), .S0 (nx1742)) ;
    xnor2 ix2372 (.Y (nx2371), .A0 (nx2373), .A1 (nx2375)) ;
    nand02_2x ix2376 (.Y (nx2375), .A0 (input_b[17]), .A1 (input_a[3])) ;
    nand02_2x ix2378 (.Y (nx2377), .A0 (input_b[16]), .A1 (input_a[5])) ;
    xnor2 ix2380 (.Y (nx2379), .A0 (nx2381), .A1 (nx2377)) ;
    xnor2 ix2382 (.Y (nx2381), .A0 (nx2383), .A1 (nx2385)) ;
    mux21_ni ix2384 (.Y (nx2383), .A0 (nx2367), .A1 (nx2375), .S0 (nx2371)) ;
    xnor2 ix2386 (.Y (nx2385), .A0 (nx2387), .A1 (nx2389)) ;
    xnor2 ix2388 (.Y (nx2387), .A0 (nx1969), .A1 (nx1989)) ;
    nand02_2x ix2390 (.Y (nx2389), .A0 (input_b[17]), .A1 (input_a[4])) ;
    xnor2 ix3231 (.Y (nx3230), .A0 (nx3226), .A1 (nx2319)) ;
    xnor2 ix3227 (.Y (nx3226), .A0 (nx2395), .A1 (nx3224)) ;
    mux21_ni ix2396 (.Y (nx2395), .A0 (nx2383), .A1 (nx2389), .S0 (nx2385)) ;
    xnor2 ix3225 (.Y (nx3224), .A0 (nx3220), .A1 (nx2401)) ;
    xnor2 ix3221 (.Y (nx3220), .A0 (nx1967), .A1 (nx3218)) ;
    nand02_2x ix2402 (.Y (nx2401), .A0 (input_b[17]), .A1 (input_a[5])) ;
    xnor2 ix3829 (.Y (nx3828), .A0 (nx3824), .A1 (nx2315)) ;
    xnor2 ix3825 (.Y (nx3824), .A0 (nx2407), .A1 (nx3822)) ;
    mux21_ni ix2408 (.Y (nx2407), .A0 (nx2401), .A1 (nx2395), .S0 (nx3224)) ;
    xnor2 ix3823 (.Y (nx3822), .A0 (nx3818), .A1 (nx2413)) ;
    xnor2 ix3819 (.Y (nx3818), .A0 (nx1963), .A1 (nx3816)) ;
    nand02_2x ix2414 (.Y (nx2413), .A0 (input_b[17]), .A1 (input_a[6])) ;
    nand02_2x ix2416 (.Y (nx2415), .A0 (input_b[16]), .A1 (input_a[8])) ;
    xnor2 ix2418 (.Y (nx2417), .A0 (nx2419), .A1 (nx2415)) ;
    xnor2 ix2420 (.Y (nx2419), .A0 (nx2421), .A1 (nx2423)) ;
    mux21_ni ix2422 (.Y (nx2421), .A0 (nx2413), .A1 (nx2407), .S0 (nx3822)) ;
    xnor2 ix2424 (.Y (nx2423), .A0 (nx2425), .A1 (nx2427)) ;
    xnor2 ix2426 (.Y (nx2425), .A0 (nx1959), .A1 (nx2031)) ;
    nand02_2x ix2428 (.Y (nx2427), .A0 (input_b[17]), .A1 (input_a[7])) ;
    xnor2 ix5835 (.Y (nx5834), .A0 (nx5832), .A1 (nx2309)) ;
    xnor2 ix5833 (.Y (nx5832), .A0 (nx2433), .A1 (nx5592)) ;
    mux21_ni ix2434 (.Y (nx2433), .A0 (nx2421), .A1 (nx2427), .S0 (nx2423)) ;
    xnor2 ix5593 (.Y (nx5592), .A0 (nx5590), .A1 (nx2439)) ;
    xnor2 ix5591 (.Y (nx5590), .A0 (nx1957), .A1 (nx5336)) ;
    nand02_2x ix2440 (.Y (nx2439), .A0 (input_b[17]), .A1 (input_a[8])) ;
    nand02_2x ix2442 (.Y (nx2441), .A0 (input_b[16]), .A1 (input_a[10])) ;
    xnor2 ix2444 (.Y (nx2443), .A0 (nx2445), .A1 (nx2441)) ;
    xnor2 ix2446 (.Y (nx2445), .A0 (nx2447), .A1 (nx2449)) ;
    mux21_ni ix2448 (.Y (nx2447), .A0 (nx2439), .A1 (nx2433), .S0 (nx5592)) ;
    xnor2 ix2450 (.Y (nx2449), .A0 (nx2451), .A1 (nx2453)) ;
    xnor2 ix2452 (.Y (nx2451), .A0 (nx1953), .A1 (nx2057)) ;
    nand02_2x ix2454 (.Y (nx2453), .A0 (input_b[17]), .A1 (input_a[9])) ;
    xnor2 ix5815 (.Y (nx5814), .A0 (nx5812), .A1 (nx2303)) ;
    xnor2 ix5813 (.Y (nx5812), .A0 (nx2459), .A1 (nx5572)) ;
    mux21_ni ix2460 (.Y (nx2459), .A0 (nx2447), .A1 (nx2453), .S0 (nx2449)) ;
    xnor2 ix5573 (.Y (nx5572), .A0 (nx5570), .A1 (nx2465)) ;
    xnor2 ix5571 (.Y (nx5570), .A0 (nx1951), .A1 (nx5316)) ;
    nand02_2x ix2466 (.Y (nx2465), .A0 (input_b[17]), .A1 (input_a[10])) ;
    nand02_2x ix2468 (.Y (nx2467), .A0 (input_b[16]), .A1 (input_a[12])) ;
    xnor2 ix2470 (.Y (nx2469), .A0 (nx2471), .A1 (nx2467)) ;
    xnor2 ix2472 (.Y (nx2471), .A0 (nx2473), .A1 (nx2475)) ;
    mux21_ni ix2474 (.Y (nx2473), .A0 (nx2465), .A1 (nx2459), .S0 (nx5572)) ;
    xnor2 ix2476 (.Y (nx2475), .A0 (nx2477), .A1 (nx2479)) ;
    xnor2 ix2478 (.Y (nx2477), .A0 (nx1947), .A1 (nx2083)) ;
    nand02_2x ix2480 (.Y (nx2479), .A0 (input_b[17]), .A1 (input_a[11])) ;
    xnor2 ix5795 (.Y (nx5794), .A0 (nx5792), .A1 (nx2297)) ;
    xnor2 ix5793 (.Y (nx5792), .A0 (nx2485), .A1 (nx5552)) ;
    mux21_ni ix2486 (.Y (nx2485), .A0 (nx2473), .A1 (nx2479), .S0 (nx2475)) ;
    xnor2 ix5553 (.Y (nx5552), .A0 (nx5550), .A1 (nx2491)) ;
    xnor2 ix5551 (.Y (nx5550), .A0 (nx1945), .A1 (nx5296)) ;
    nand02_2x ix2492 (.Y (nx2491), .A0 (input_b[17]), .A1 (input_a[12])) ;
    nand02_2x ix2494 (.Y (nx2493), .A0 (input_b[16]), .A1 (input_a[14])) ;
    xnor2 ix2496 (.Y (nx2495), .A0 (nx2497), .A1 (nx2493)) ;
    xnor2 ix2498 (.Y (nx2497), .A0 (nx2499), .A1 (nx2501)) ;
    mux21_ni ix2500 (.Y (nx2499), .A0 (nx2491), .A1 (nx2485), .S0 (nx5552)) ;
    xnor2 ix2502 (.Y (nx2501), .A0 (nx2503), .A1 (nx2505)) ;
    xnor2 ix2504 (.Y (nx2503), .A0 (nx1941), .A1 (nx2109)) ;
    nand02_2x ix2506 (.Y (nx2505), .A0 (input_b[17]), .A1 (input_a[13])) ;
    xnor2 ix5775 (.Y (nx5774), .A0 (nx5772), .A1 (nx2291)) ;
    xnor2 ix5773 (.Y (nx5772), .A0 (nx2511), .A1 (nx5532)) ;
    mux21_ni ix2512 (.Y (nx2511), .A0 (nx2499), .A1 (nx2505), .S0 (nx2501)) ;
    xnor2 ix5533 (.Y (nx5532), .A0 (nx5530), .A1 (nx2517)) ;
    xnor2 ix5531 (.Y (nx5530), .A0 (nx1939), .A1 (nx5276)) ;
    nand02_2x ix2518 (.Y (nx2517), .A0 (input_b[17]), .A1 (input_a[14])) ;
    nand02_2x ix2520 (.Y (nx2519), .A0 (input_b[16]), .A1 (input_a[16])) ;
    xnor2 ix2522 (.Y (nx2521), .A0 (nx2523), .A1 (nx2519)) ;
    xnor2 ix2524 (.Y (nx2523), .A0 (nx2525), .A1 (nx2527)) ;
    mux21_ni ix2526 (.Y (nx2525), .A0 (nx2517), .A1 (nx2511), .S0 (nx5532)) ;
    xnor2 ix2528 (.Y (nx2527), .A0 (nx2529), .A1 (nx2531)) ;
    xnor2 ix2530 (.Y (nx2529), .A0 (nx1935), .A1 (nx2135)) ;
    nand02_2x ix2532 (.Y (nx2531), .A0 (input_b[17]), .A1 (input_a[15])) ;
    xnor2 ix5755 (.Y (nx5754), .A0 (nx5752), .A1 (nx2285)) ;
    xnor2 ix5753 (.Y (nx5752), .A0 (nx2537), .A1 (nx5512)) ;
    mux21_ni ix2538 (.Y (nx2537), .A0 (nx2525), .A1 (nx2531), .S0 (nx2527)) ;
    xnor2 ix5513 (.Y (nx5512), .A0 (nx5510), .A1 (nx2543)) ;
    xnor2 ix5511 (.Y (nx5510), .A0 (nx1933), .A1 (nx5256)) ;
    nand02_2x ix2544 (.Y (nx2543), .A0 (input_b[17]), .A1 (input_a[16])) ;
    nand02_2x ix2546 (.Y (nx2545), .A0 (input_b[16]), .A1 (input_a[18])) ;
    xnor2 ix2548 (.Y (nx2547), .A0 (nx2549), .A1 (nx2545)) ;
    xnor2 ix2550 (.Y (nx2549), .A0 (nx2551), .A1 (nx2553)) ;
    mux21_ni ix2552 (.Y (nx2551), .A0 (nx2543), .A1 (nx2537), .S0 (nx5512)) ;
    xnor2 ix2554 (.Y (nx2553), .A0 (nx2555), .A1 (nx2557)) ;
    xnor2 ix2556 (.Y (nx2555), .A0 (nx1929), .A1 (nx2161)) ;
    nand02_2x ix2558 (.Y (nx2557), .A0 (input_b[17]), .A1 (input_a[17])) ;
    xnor2 ix5735 (.Y (nx5734), .A0 (nx5732), .A1 (nx2279)) ;
    xnor2 ix5733 (.Y (nx5732), .A0 (nx2563), .A1 (nx5492)) ;
    mux21_ni ix2564 (.Y (nx2563), .A0 (nx2551), .A1 (nx2557), .S0 (nx2553)) ;
    xnor2 ix5493 (.Y (nx5492), .A0 (nx5490), .A1 (nx2569)) ;
    xnor2 ix5491 (.Y (nx5490), .A0 (nx1927), .A1 (nx5236)) ;
    nand02_2x ix2570 (.Y (nx2569), .A0 (input_b[17]), .A1 (input_a[18])) ;
    nand02_2x ix2572 (.Y (nx2571), .A0 (input_b[16]), .A1 (input_a[20])) ;
    xnor2 ix2574 (.Y (nx2573), .A0 (nx2575), .A1 (nx2571)) ;
    xnor2 ix2576 (.Y (nx2575), .A0 (nx2577), .A1 (nx2579)) ;
    mux21_ni ix2578 (.Y (nx2577), .A0 (nx2569), .A1 (nx2563), .S0 (nx5492)) ;
    xnor2 ix2580 (.Y (nx2579), .A0 (nx2581), .A1 (nx2583)) ;
    xnor2 ix2582 (.Y (nx2581), .A0 (nx1923), .A1 (nx2187)) ;
    nand02_2x ix2584 (.Y (nx2583), .A0 (input_b[17]), .A1 (input_a[19])) ;
    xnor2 ix5715 (.Y (nx5714), .A0 (nx5712), .A1 (nx2273)) ;
    xnor2 ix5713 (.Y (nx5712), .A0 (nx2589), .A1 (nx5472)) ;
    mux21_ni ix2590 (.Y (nx2589), .A0 (nx2577), .A1 (nx2583), .S0 (nx2579)) ;
    xnor2 ix5473 (.Y (nx5472), .A0 (nx5470), .A1 (nx2595)) ;
    xnor2 ix5471 (.Y (nx5470), .A0 (nx1921), .A1 (nx5216)) ;
    nand02_2x ix2596 (.Y (nx2595), .A0 (input_b[17]), .A1 (input_a[20])) ;
    nand02_2x ix2598 (.Y (nx2597), .A0 (input_b[16]), .A1 (input_a[22])) ;
    xnor2 ix2600 (.Y (nx2599), .A0 (nx2601), .A1 (nx2597)) ;
    xnor2 ix2602 (.Y (nx2601), .A0 (nx2603), .A1 (nx2605)) ;
    mux21_ni ix2604 (.Y (nx2603), .A0 (nx2595), .A1 (nx2589), .S0 (nx5472)) ;
    xnor2 ix2606 (.Y (nx2605), .A0 (nx2607), .A1 (nx2609)) ;
    xnor2 ix2608 (.Y (nx2607), .A0 (nx1917), .A1 (nx2213)) ;
    nand02_2x ix2610 (.Y (nx2609), .A0 (input_b[17]), .A1 (input_a[21])) ;
    xnor2 ix2612 (.Y (nx2611), .A0 (input_b[16]), .A1 (nx5692)) ;
    xnor2 ix5693 (.Y (nx5692), .A0 (nx2615), .A1 (nx5452)) ;
    mux21_ni ix2616 (.Y (nx2615), .A0 (nx2603), .A1 (nx2609), .S0 (nx2605)) ;
    xnor2 ix5453 (.Y (nx5452), .A0 (nx5450), .A1 (nx2621)) ;
    xnor2 ix5451 (.Y (nx5450), .A0 (nx1915), .A1 (nx5196)) ;
    nand02_2x ix2622 (.Y (nx2621), .A0 (input_b[17]), .A1 (input_a[22])) ;
    mux21_ni ix7885 (.Y (nx7884), .A0 (nx7880), .A1 (nx6152), .S0 (nx5655)) ;
    xnor2 ix2628 (.Y (nx2627), .A0 (nx2629), .A1 (nx2971)) ;
    mux21_ni ix2630 (.Y (nx2629), .A0 (nx2631), .A1 (nx2957), .S0 (nx2959)) ;
    mux21_ni ix2632 (.Y (nx2631), .A0 (nx2633), .A1 (nx2635), .S0 (nx6176)) ;
    nand02_2x ix2634 (.Y (nx2633), .A0 (input_b[14]), .A1 (input_a[21])) ;
    mux21_ni ix2636 (.Y (nx2635), .A0 (nx2637), .A1 (nx2931), .S0 (nx2933)) ;
    mux21_ni ix2638 (.Y (nx2637), .A0 (nx2639), .A1 (nx2641), .S0 (nx6196)) ;
    nand02_2x ix2640 (.Y (nx2639), .A0 (input_b[14]), .A1 (input_a[19])) ;
    mux21_ni ix2642 (.Y (nx2641), .A0 (nx2643), .A1 (nx2905), .S0 (nx2907)) ;
    mux21_ni ix2644 (.Y (nx2643), .A0 (nx2645), .A1 (nx2647), .S0 (nx6216)) ;
    nand02_2x ix2646 (.Y (nx2645), .A0 (input_b[14]), .A1 (input_a[17])) ;
    mux21_ni ix2648 (.Y (nx2647), .A0 (nx2649), .A1 (nx2879), .S0 (nx2881)) ;
    mux21_ni ix2650 (.Y (nx2649), .A0 (nx2651), .A1 (nx2653), .S0 (nx6236)) ;
    nand02_2x ix2652 (.Y (nx2651), .A0 (input_b[14]), .A1 (input_a[15])) ;
    mux21_ni ix2654 (.Y (nx2653), .A0 (nx2655), .A1 (nx2853), .S0 (nx2855)) ;
    mux21_ni ix2656 (.Y (nx2655), .A0 (nx2657), .A1 (nx2659), .S0 (nx6256)) ;
    nand02_2x ix2658 (.Y (nx2657), .A0 (input_b[14]), .A1 (input_a[13])) ;
    mux21_ni ix2660 (.Y (nx2659), .A0 (nx2661), .A1 (nx2827), .S0 (nx2829)) ;
    mux21_ni ix2662 (.Y (nx2661), .A0 (nx2663), .A1 (nx2665), .S0 (nx6276)) ;
    nand02_2x ix2664 (.Y (nx2663), .A0 (input_b[14]), .A1 (input_a[11])) ;
    mux21_ni ix2666 (.Y (nx2665), .A0 (nx2667), .A1 (nx2801), .S0 (nx2803)) ;
    mux21_ni ix2668 (.Y (nx2667), .A0 (nx2669), .A1 (nx2671), .S0 (nx3840)) ;
    nand02_2x ix2670 (.Y (nx2669), .A0 (input_b[14]), .A1 (input_a[9])) ;
    mux21_ni ix2672 (.Y (nx2671), .A0 (nx2673), .A1 (nx2675), .S0 (nx3242)) ;
    nand02_2x ix2674 (.Y (nx2673), .A0 (input_b[14]), .A1 (input_a[8])) ;
    mux21_ni ix2676 (.Y (nx2675), .A0 (nx2677), .A1 (nx2763), .S0 (nx2765)) ;
    mux21_ni ix2678 (.Y (nx2677), .A0 (nx2679), .A1 (nx2749), .S0 (nx2751)) ;
    mux21_ni ix2680 (.Y (nx2679), .A0 (nx2681), .A1 (nx2735), .S0 (nx2737)) ;
    mux21_ni ix2682 (.Y (nx2681), .A0 (nx2683), .A1 (nx2719), .S0 (nx2721)) ;
    mux21_ni ix2684 (.Y (nx2683), .A0 (nx2685), .A1 (nx2703), .S0 (nx2705)) ;
    mux21_ni ix2686 (.Y (nx2685), .A0 (nx2687), .A1 (nx2689), .S0 (nx782)) ;
    nand02_2x ix2688 (.Y (nx2687), .A0 (input_b[14]), .A1 (input_a[2])) ;
    xnor2 ix783 (.Y (nx782), .A0 (nx778), .A1 (nx2687)) ;
    inv02 ix2698 (.Y (nx2697), .A (input_b[15])) ;
    inv02 ix2700 (.Y (nx2699), .A (input_b[16])) ;
    aoi22 ix2702 (.Y (nx2701), .A0 (input_b[16]), .A1 (input_a[0]), .B0 (
          input_b[15]), .B1 (input_a[1])) ;
    nand02_2x ix2704 (.Y (nx2703), .A0 (input_b[14]), .A1 (input_a[3])) ;
    xnor2 ix2706 (.Y (nx2705), .A0 (nx2707), .A1 (nx2703)) ;
    xnor2 ix1047 (.Y (nx1046), .A0 (nx1042), .A1 (nx2717)) ;
    aoi22 ix2716 (.Y (nx2715), .A0 (input_b[17]), .A1 (input_a[0]), .B0 (
          input_b[16]), .B1 (input_a[1])) ;
    nand02_2x ix2718 (.Y (nx2717), .A0 (input_b[15]), .A1 (input_a[2])) ;
    nand02_2x ix2720 (.Y (nx2719), .A0 (input_b[14]), .A1 (input_a[4])) ;
    xnor2 ix2722 (.Y (nx2721), .A0 (nx2723), .A1 (nx2719)) ;
    xnor2 ix2724 (.Y (nx2723), .A0 (nx2725), .A1 (nx2729)) ;
    mux21_ni ix2726 (.Y (nx2725), .A0 (nx2717), .A1 (nx2727), .S0 (nx1046)) ;
    xnor2 ix2730 (.Y (nx2729), .A0 (nx2731), .A1 (nx2733)) ;
    nand02_2x ix2734 (.Y (nx2733), .A0 (input_b[15]), .A1 (input_a[3])) ;
    nand02_2x ix2736 (.Y (nx2735), .A0 (input_b[14]), .A1 (input_a[5])) ;
    xnor2 ix2738 (.Y (nx2737), .A0 (nx2739), .A1 (nx2735)) ;
    xnor2 ix2740 (.Y (nx2739), .A0 (nx2741), .A1 (nx2743)) ;
    mux21_ni ix2742 (.Y (nx2741), .A0 (nx2725), .A1 (nx2733), .S0 (nx2729)) ;
    xnor2 ix2744 (.Y (nx2743), .A0 (nx2745), .A1 (nx2747)) ;
    xnor2 ix2746 (.Y (nx2745), .A0 (nx2327), .A1 (nx2347)) ;
    nand02_2x ix2748 (.Y (nx2747), .A0 (input_b[15]), .A1 (input_a[4])) ;
    nand02_2x ix2750 (.Y (nx2749), .A0 (input_b[14]), .A1 (input_a[6])) ;
    xnor2 ix2752 (.Y (nx2751), .A0 (nx2753), .A1 (nx2749)) ;
    xnor2 ix2754 (.Y (nx2753), .A0 (nx2755), .A1 (nx2757)) ;
    mux21_ni ix2756 (.Y (nx2755), .A0 (nx2741), .A1 (nx2747), .S0 (nx2743)) ;
    xnor2 ix2758 (.Y (nx2757), .A0 (nx2759), .A1 (nx2761)) ;
    xnor2 ix2760 (.Y (nx2759), .A0 (nx2325), .A1 (nx2363)) ;
    nand02_2x ix2762 (.Y (nx2761), .A0 (input_b[15]), .A1 (input_a[5])) ;
    nand02_2x ix2764 (.Y (nx2763), .A0 (input_b[14]), .A1 (input_a[7])) ;
    xnor2 ix2766 (.Y (nx2765), .A0 (nx2767), .A1 (nx2763)) ;
    xnor2 ix2768 (.Y (nx2767), .A0 (nx2769), .A1 (nx2771)) ;
    mux21_ni ix2770 (.Y (nx2769), .A0 (nx2755), .A1 (nx2761), .S0 (nx2757)) ;
    xnor2 ix2772 (.Y (nx2771), .A0 (nx2773), .A1 (nx2775)) ;
    xnor2 ix2774 (.Y (nx2773), .A0 (nx2323), .A1 (nx2379)) ;
    nand02_2x ix2776 (.Y (nx2775), .A0 (input_b[15]), .A1 (input_a[6])) ;
    xnor2 ix3243 (.Y (nx3242), .A0 (nx3238), .A1 (nx2673)) ;
    xnor2 ix3239 (.Y (nx3238), .A0 (nx2781), .A1 (nx3236)) ;
    mux21_ni ix2782 (.Y (nx2781), .A0 (nx2769), .A1 (nx2775), .S0 (nx2771)) ;
    xnor2 ix3237 (.Y (nx3236), .A0 (nx3232), .A1 (nx2787)) ;
    xnor2 ix3233 (.Y (nx3232), .A0 (nx2321), .A1 (nx3230)) ;
    nand02_2x ix2788 (.Y (nx2787), .A0 (input_b[15]), .A1 (input_a[7])) ;
    xnor2 ix3841 (.Y (nx3840), .A0 (nx3836), .A1 (nx2669)) ;
    xnor2 ix3837 (.Y (nx3836), .A0 (nx2793), .A1 (nx3834)) ;
    mux21_ni ix2794 (.Y (nx2793), .A0 (nx2787), .A1 (nx2781), .S0 (nx3236)) ;
    xnor2 ix3835 (.Y (nx3834), .A0 (nx3830), .A1 (nx2799)) ;
    xnor2 ix3831 (.Y (nx3830), .A0 (nx2317), .A1 (nx3828)) ;
    nand02_2x ix2800 (.Y (nx2799), .A0 (input_b[15]), .A1 (input_a[8])) ;
    nand02_2x ix2802 (.Y (nx2801), .A0 (input_b[14]), .A1 (input_a[10])) ;
    xnor2 ix2804 (.Y (nx2803), .A0 (nx2805), .A1 (nx2801)) ;
    xnor2 ix2806 (.Y (nx2805), .A0 (nx2807), .A1 (nx2809)) ;
    mux21_ni ix2808 (.Y (nx2807), .A0 (nx2799), .A1 (nx2793), .S0 (nx3834)) ;
    xnor2 ix2810 (.Y (nx2809), .A0 (nx2811), .A1 (nx2813)) ;
    xnor2 ix2812 (.Y (nx2811), .A0 (nx2313), .A1 (nx2417)) ;
    nand02_2x ix2814 (.Y (nx2813), .A0 (input_b[15]), .A1 (input_a[9])) ;
    xnor2 ix6277 (.Y (nx6276), .A0 (nx6274), .A1 (nx2663)) ;
    xnor2 ix6275 (.Y (nx6274), .A0 (nx2819), .A1 (nx6062)) ;
    mux21_ni ix2820 (.Y (nx2819), .A0 (nx2807), .A1 (nx2813), .S0 (nx2809)) ;
    xnor2 ix6063 (.Y (nx6062), .A0 (nx6060), .A1 (nx2825)) ;
    xnor2 ix6061 (.Y (nx6060), .A0 (nx2311), .A1 (nx5834)) ;
    nand02_2x ix2826 (.Y (nx2825), .A0 (input_b[15]), .A1 (input_a[10])) ;
    nand02_2x ix2828 (.Y (nx2827), .A0 (input_b[14]), .A1 (input_a[12])) ;
    xnor2 ix2830 (.Y (nx2829), .A0 (nx2831), .A1 (nx2827)) ;
    xnor2 ix2832 (.Y (nx2831), .A0 (nx2833), .A1 (nx2835)) ;
    mux21_ni ix2834 (.Y (nx2833), .A0 (nx2825), .A1 (nx2819), .S0 (nx6062)) ;
    xnor2 ix2836 (.Y (nx2835), .A0 (nx2837), .A1 (nx2839)) ;
    xnor2 ix2838 (.Y (nx2837), .A0 (nx2307), .A1 (nx2443)) ;
    nand02_2x ix2840 (.Y (nx2839), .A0 (input_b[15]), .A1 (input_a[11])) ;
    xnor2 ix6257 (.Y (nx6256), .A0 (nx6254), .A1 (nx2657)) ;
    xnor2 ix6255 (.Y (nx6254), .A0 (nx2845), .A1 (nx6042)) ;
    mux21_ni ix2846 (.Y (nx2845), .A0 (nx2833), .A1 (nx2839), .S0 (nx2835)) ;
    xnor2 ix6043 (.Y (nx6042), .A0 (nx6040), .A1 (nx2851)) ;
    xnor2 ix6041 (.Y (nx6040), .A0 (nx2305), .A1 (nx5814)) ;
    nand02_2x ix2852 (.Y (nx2851), .A0 (input_b[15]), .A1 (input_a[12])) ;
    nand02_2x ix2854 (.Y (nx2853), .A0 (input_b[14]), .A1 (input_a[14])) ;
    xnor2 ix2856 (.Y (nx2855), .A0 (nx2857), .A1 (nx2853)) ;
    xnor2 ix2858 (.Y (nx2857), .A0 (nx2859), .A1 (nx2861)) ;
    mux21_ni ix2860 (.Y (nx2859), .A0 (nx2851), .A1 (nx2845), .S0 (nx6042)) ;
    xnor2 ix2862 (.Y (nx2861), .A0 (nx2863), .A1 (nx2865)) ;
    xnor2 ix2864 (.Y (nx2863), .A0 (nx2301), .A1 (nx2469)) ;
    nand02_2x ix2866 (.Y (nx2865), .A0 (input_b[15]), .A1 (input_a[13])) ;
    xnor2 ix6237 (.Y (nx6236), .A0 (nx6234), .A1 (nx2651)) ;
    xnor2 ix6235 (.Y (nx6234), .A0 (nx2871), .A1 (nx6022)) ;
    mux21_ni ix2872 (.Y (nx2871), .A0 (nx2859), .A1 (nx2865), .S0 (nx2861)) ;
    xnor2 ix6023 (.Y (nx6022), .A0 (nx6020), .A1 (nx2877)) ;
    xnor2 ix6021 (.Y (nx6020), .A0 (nx2299), .A1 (nx5794)) ;
    nand02_2x ix2878 (.Y (nx2877), .A0 (input_b[15]), .A1 (input_a[14])) ;
    nand02_2x ix2880 (.Y (nx2879), .A0 (input_b[14]), .A1 (input_a[16])) ;
    xnor2 ix2882 (.Y (nx2881), .A0 (nx2883), .A1 (nx2879)) ;
    xnor2 ix2884 (.Y (nx2883), .A0 (nx2885), .A1 (nx2887)) ;
    mux21_ni ix2886 (.Y (nx2885), .A0 (nx2877), .A1 (nx2871), .S0 (nx6022)) ;
    xnor2 ix2888 (.Y (nx2887), .A0 (nx2889), .A1 (nx2891)) ;
    xnor2 ix2890 (.Y (nx2889), .A0 (nx2295), .A1 (nx2495)) ;
    nand02_2x ix2892 (.Y (nx2891), .A0 (input_b[15]), .A1 (input_a[15])) ;
    xnor2 ix6217 (.Y (nx6216), .A0 (nx6214), .A1 (nx2645)) ;
    xnor2 ix6215 (.Y (nx6214), .A0 (nx2897), .A1 (nx6002)) ;
    mux21_ni ix2898 (.Y (nx2897), .A0 (nx2885), .A1 (nx2891), .S0 (nx2887)) ;
    xnor2 ix6003 (.Y (nx6002), .A0 (nx6000), .A1 (nx2903)) ;
    xnor2 ix6001 (.Y (nx6000), .A0 (nx2293), .A1 (nx5774)) ;
    nand02_2x ix2904 (.Y (nx2903), .A0 (input_b[15]), .A1 (input_a[16])) ;
    nand02_2x ix2906 (.Y (nx2905), .A0 (input_b[14]), .A1 (input_a[18])) ;
    xnor2 ix2908 (.Y (nx2907), .A0 (nx2909), .A1 (nx2905)) ;
    xnor2 ix2910 (.Y (nx2909), .A0 (nx2911), .A1 (nx2913)) ;
    mux21_ni ix2912 (.Y (nx2911), .A0 (nx2903), .A1 (nx2897), .S0 (nx6002)) ;
    xnor2 ix2914 (.Y (nx2913), .A0 (nx2915), .A1 (nx2917)) ;
    xnor2 ix2916 (.Y (nx2915), .A0 (nx2289), .A1 (nx2521)) ;
    nand02_2x ix2918 (.Y (nx2917), .A0 (input_b[15]), .A1 (input_a[17])) ;
    xnor2 ix6197 (.Y (nx6196), .A0 (nx6194), .A1 (nx2639)) ;
    xnor2 ix6195 (.Y (nx6194), .A0 (nx2923), .A1 (nx5982)) ;
    mux21_ni ix2924 (.Y (nx2923), .A0 (nx2911), .A1 (nx2917), .S0 (nx2913)) ;
    xnor2 ix5983 (.Y (nx5982), .A0 (nx5980), .A1 (nx2929)) ;
    xnor2 ix5981 (.Y (nx5980), .A0 (nx2287), .A1 (nx5754)) ;
    nand02_2x ix2930 (.Y (nx2929), .A0 (input_b[15]), .A1 (input_a[18])) ;
    nand02_2x ix2932 (.Y (nx2931), .A0 (input_b[14]), .A1 (input_a[20])) ;
    xnor2 ix2934 (.Y (nx2933), .A0 (nx2935), .A1 (nx2931)) ;
    xnor2 ix2936 (.Y (nx2935), .A0 (nx2937), .A1 (nx2939)) ;
    mux21_ni ix2938 (.Y (nx2937), .A0 (nx2929), .A1 (nx2923), .S0 (nx5982)) ;
    xnor2 ix2940 (.Y (nx2939), .A0 (nx2941), .A1 (nx2943)) ;
    xnor2 ix2942 (.Y (nx2941), .A0 (nx2283), .A1 (nx2547)) ;
    nand02_2x ix2944 (.Y (nx2943), .A0 (input_b[15]), .A1 (input_a[19])) ;
    xnor2 ix6177 (.Y (nx6176), .A0 (nx6174), .A1 (nx2633)) ;
    xnor2 ix6175 (.Y (nx6174), .A0 (nx2949), .A1 (nx5962)) ;
    mux21_ni ix2950 (.Y (nx2949), .A0 (nx2937), .A1 (nx2943), .S0 (nx2939)) ;
    xnor2 ix5963 (.Y (nx5962), .A0 (nx5960), .A1 (nx2955)) ;
    xnor2 ix5961 (.Y (nx5960), .A0 (nx2281), .A1 (nx5734)) ;
    nand02_2x ix2956 (.Y (nx2955), .A0 (input_b[15]), .A1 (input_a[20])) ;
    nand02_2x ix2958 (.Y (nx2957), .A0 (input_b[14]), .A1 (input_a[22])) ;
    xnor2 ix2960 (.Y (nx2959), .A0 (nx2961), .A1 (nx2957)) ;
    xnor2 ix2962 (.Y (nx2961), .A0 (nx2963), .A1 (nx2965)) ;
    mux21_ni ix2964 (.Y (nx2963), .A0 (nx2955), .A1 (nx2949), .S0 (nx5962)) ;
    xnor2 ix2966 (.Y (nx2965), .A0 (nx2967), .A1 (nx2969)) ;
    xnor2 ix2968 (.Y (nx2967), .A0 (nx2277), .A1 (nx2573)) ;
    nand02_2x ix2970 (.Y (nx2969), .A0 (input_b[15]), .A1 (input_a[21])) ;
    xnor2 ix2972 (.Y (nx2971), .A0 (input_b[14]), .A1 (nx6154)) ;
    xnor2 ix6155 (.Y (nx6154), .A0 (nx2975), .A1 (nx5942)) ;
    mux21_ni ix2976 (.Y (nx2975), .A0 (nx2963), .A1 (nx2969), .S0 (nx2965)) ;
    xnor2 ix5943 (.Y (nx5942), .A0 (nx5940), .A1 (nx2981)) ;
    xnor2 ix5941 (.Y (nx5940), .A0 (nx2275), .A1 (nx5714)) ;
    nand02_2x ix2982 (.Y (nx2981), .A0 (input_b[15]), .A1 (input_a[22])) ;
    mux21_ni ix2984 (.Y (nx2983), .A0 (nx2985), .A1 (nx5625), .S0 (nx5633)) ;
    mux21_ni ix2986 (.Y (nx2985), .A0 (nx2987), .A1 (nx3343), .S0 (nx6902)) ;
    xnor2 ix2988 (.Y (nx2987), .A0 (nx2989), .A1 (nx3331)) ;
    mux21_ni ix2990 (.Y (nx2989), .A0 (nx2991), .A1 (nx3317), .S0 (nx3319)) ;
    mux21_ni ix2992 (.Y (nx2991), .A0 (nx2993), .A1 (nx2995), .S0 (nx6582)) ;
    nand02_2x ix2994 (.Y (nx2993), .A0 (input_b[12]), .A1 (input_a[21])) ;
    mux21_ni ix2996 (.Y (nx2995), .A0 (nx2997), .A1 (nx3291), .S0 (nx3293)) ;
    mux21_ni ix2998 (.Y (nx2997), .A0 (nx2999), .A1 (nx3001), .S0 (nx6602)) ;
    nand02_2x ix3000 (.Y (nx2999), .A0 (input_b[12]), .A1 (input_a[19])) ;
    mux21_ni ix3002 (.Y (nx3001), .A0 (nx3003), .A1 (nx3265), .S0 (nx3267)) ;
    mux21_ni ix3004 (.Y (nx3003), .A0 (nx3005), .A1 (nx3007), .S0 (nx6622)) ;
    nand02_2x ix3006 (.Y (nx3005), .A0 (input_b[12]), .A1 (input_a[17])) ;
    mux21_ni ix3008 (.Y (nx3007), .A0 (nx3009), .A1 (nx3239), .S0 (nx3241)) ;
    mux21_ni ix3010 (.Y (nx3009), .A0 (nx3011), .A1 (nx3013), .S0 (nx6642)) ;
    nand02_2x ix3012 (.Y (nx3011), .A0 (input_b[12]), .A1 (input_a[15])) ;
    mux21_ni ix3014 (.Y (nx3013), .A0 (nx3015), .A1 (nx3213), .S0 (nx3215)) ;
    mux21_ni ix3016 (.Y (nx3015), .A0 (nx3017), .A1 (nx3019), .S0 (nx6662)) ;
    nand02_2x ix3018 (.Y (nx3017), .A0 (input_b[12]), .A1 (input_a[13])) ;
    mux21_ni ix3020 (.Y (nx3019), .A0 (nx3021), .A1 (nx3187), .S0 (nx3189)) ;
    mux21_ni ix3022 (.Y (nx3021), .A0 (nx3023), .A1 (nx3025), .S0 (nx3852)) ;
    nand02_2x ix3024 (.Y (nx3023), .A0 (input_b[12]), .A1 (input_a[11])) ;
    mux21_ni ix3026 (.Y (nx3025), .A0 (nx3027), .A1 (nx3029), .S0 (nx3254)) ;
    nand02_2x ix3028 (.Y (nx3027), .A0 (input_b[12]), .A1 (input_a[10])) ;
    mux21_ni ix3030 (.Y (nx3029), .A0 (nx3031), .A1 (nx3149), .S0 (nx3151)) ;
    mux21_ni ix3032 (.Y (nx3031), .A0 (nx3033), .A1 (nx3135), .S0 (nx3137)) ;
    mux21_ni ix3034 (.Y (nx3033), .A0 (nx3035), .A1 (nx3121), .S0 (nx3123)) ;
    mux21_ni ix3036 (.Y (nx3035), .A0 (nx3037), .A1 (nx3107), .S0 (nx3109)) ;
    mux21_ni ix3038 (.Y (nx3037), .A0 (nx3039), .A1 (nx3093), .S0 (nx3095)) ;
    mux21_ni ix3040 (.Y (nx3039), .A0 (nx3041), .A1 (nx3077), .S0 (nx3079)) ;
    mux21_ni ix3042 (.Y (nx3041), .A0 (nx3043), .A1 (nx3061), .S0 (nx3063)) ;
    mux21_ni ix3044 (.Y (nx3043), .A0 (nx3045), .A1 (nx3047), .S0 (nx422)) ;
    nand02_2x ix3046 (.Y (nx3045), .A0 (input_b[12]), .A1 (input_a[2])) ;
    xnor2 ix423 (.Y (nx422), .A0 (nx418), .A1 (nx3045)) ;
    inv02 ix3056 (.Y (nx3055), .A (input_b[13])) ;
    inv02 ix3058 (.Y (nx3057), .A (input_b[14])) ;
    aoi22 ix3060 (.Y (nx3059), .A0 (input_b[14]), .A1 (input_a[0]), .B0 (
          input_b[13]), .B1 (input_a[1])) ;
    nand02_2x ix3062 (.Y (nx3061), .A0 (input_b[12]), .A1 (input_a[3])) ;
    xnor2 ix3064 (.Y (nx3063), .A0 (nx3065), .A1 (nx3061)) ;
    xnor2 ix575 (.Y (nx574), .A0 (nx570), .A1 (nx3075)) ;
    aoi22 ix3074 (.Y (nx3073), .A0 (input_b[15]), .A1 (input_a[0]), .B0 (
          input_b[14]), .B1 (input_a[1])) ;
    nand02_2x ix3076 (.Y (nx3075), .A0 (input_b[13]), .A1 (input_a[2])) ;
    nand02_2x ix3078 (.Y (nx3077), .A0 (input_b[12]), .A1 (input_a[4])) ;
    xnor2 ix3080 (.Y (nx3079), .A0 (nx3081), .A1 (nx3077)) ;
    xnor2 ix3082 (.Y (nx3081), .A0 (nx3083), .A1 (nx3087)) ;
    mux21_ni ix3084 (.Y (nx3083), .A0 (nx3075), .A1 (nx3085), .S0 (nx574)) ;
    xnor2 ix3088 (.Y (nx3087), .A0 (nx3089), .A1 (nx3091)) ;
    nand02_2x ix3092 (.Y (nx3091), .A0 (input_b[13]), .A1 (input_a[3])) ;
    nand02_2x ix3094 (.Y (nx3093), .A0 (input_b[12]), .A1 (input_a[5])) ;
    xnor2 ix3096 (.Y (nx3095), .A0 (nx3097), .A1 (nx3093)) ;
    xnor2 ix3098 (.Y (nx3097), .A0 (nx3099), .A1 (nx3101)) ;
    mux21_ni ix3100 (.Y (nx3099), .A0 (nx3083), .A1 (nx3091), .S0 (nx3087)) ;
    xnor2 ix3102 (.Y (nx3101), .A0 (nx3103), .A1 (nx3105)) ;
    xnor2 ix3104 (.Y (nx3103), .A0 (nx2685), .A1 (nx2705)) ;
    nand02_2x ix3106 (.Y (nx3105), .A0 (input_b[13]), .A1 (input_a[4])) ;
    nand02_2x ix3108 (.Y (nx3107), .A0 (input_b[12]), .A1 (input_a[6])) ;
    xnor2 ix3110 (.Y (nx3109), .A0 (nx3111), .A1 (nx3107)) ;
    xnor2 ix3112 (.Y (nx3111), .A0 (nx3113), .A1 (nx3115)) ;
    mux21_ni ix3114 (.Y (nx3113), .A0 (nx3099), .A1 (nx3105), .S0 (nx3101)) ;
    xnor2 ix3116 (.Y (nx3115), .A0 (nx3117), .A1 (nx3119)) ;
    xnor2 ix3118 (.Y (nx3117), .A0 (nx2683), .A1 (nx2721)) ;
    nand02_2x ix3120 (.Y (nx3119), .A0 (input_b[13]), .A1 (input_a[5])) ;
    nand02_2x ix3122 (.Y (nx3121), .A0 (input_b[12]), .A1 (input_a[7])) ;
    xnor2 ix3124 (.Y (nx3123), .A0 (nx3125), .A1 (nx3121)) ;
    xnor2 ix3126 (.Y (nx3125), .A0 (nx3127), .A1 (nx3129)) ;
    mux21_ni ix3128 (.Y (nx3127), .A0 (nx3113), .A1 (nx3119), .S0 (nx3115)) ;
    xnor2 ix3130 (.Y (nx3129), .A0 (nx3131), .A1 (nx3133)) ;
    xnor2 ix3132 (.Y (nx3131), .A0 (nx2681), .A1 (nx2737)) ;
    nand02_2x ix3134 (.Y (nx3133), .A0 (input_b[13]), .A1 (input_a[6])) ;
    nand02_2x ix3136 (.Y (nx3135), .A0 (input_b[12]), .A1 (input_a[8])) ;
    xnor2 ix3138 (.Y (nx3137), .A0 (nx3139), .A1 (nx3135)) ;
    xnor2 ix3140 (.Y (nx3139), .A0 (nx3141), .A1 (nx3143)) ;
    mux21_ni ix3142 (.Y (nx3141), .A0 (nx3127), .A1 (nx3133), .S0 (nx3129)) ;
    xnor2 ix3144 (.Y (nx3143), .A0 (nx3145), .A1 (nx3147)) ;
    xnor2 ix3146 (.Y (nx3145), .A0 (nx2679), .A1 (nx2751)) ;
    nand02_2x ix3148 (.Y (nx3147), .A0 (input_b[13]), .A1 (input_a[7])) ;
    nand02_2x ix3150 (.Y (nx3149), .A0 (input_b[12]), .A1 (input_a[9])) ;
    xnor2 ix3152 (.Y (nx3151), .A0 (nx3153), .A1 (nx3149)) ;
    xnor2 ix3154 (.Y (nx3153), .A0 (nx3155), .A1 (nx3157)) ;
    mux21_ni ix3156 (.Y (nx3155), .A0 (nx3141), .A1 (nx3147), .S0 (nx3143)) ;
    xnor2 ix3158 (.Y (nx3157), .A0 (nx3159), .A1 (nx3161)) ;
    xnor2 ix3160 (.Y (nx3159), .A0 (nx2677), .A1 (nx2765)) ;
    nand02_2x ix3162 (.Y (nx3161), .A0 (input_b[13]), .A1 (input_a[8])) ;
    xnor2 ix3255 (.Y (nx3254), .A0 (nx3250), .A1 (nx3027)) ;
    xnor2 ix3251 (.Y (nx3250), .A0 (nx3167), .A1 (nx3248)) ;
    mux21_ni ix3168 (.Y (nx3167), .A0 (nx3155), .A1 (nx3161), .S0 (nx3157)) ;
    xnor2 ix3249 (.Y (nx3248), .A0 (nx3244), .A1 (nx3173)) ;
    xnor2 ix3245 (.Y (nx3244), .A0 (nx2675), .A1 (nx3242)) ;
    nand02_2x ix3174 (.Y (nx3173), .A0 (input_b[13]), .A1 (input_a[9])) ;
    xnor2 ix3853 (.Y (nx3852), .A0 (nx3848), .A1 (nx3023)) ;
    xnor2 ix3849 (.Y (nx3848), .A0 (nx3179), .A1 (nx3846)) ;
    mux21_ni ix3180 (.Y (nx3179), .A0 (nx3173), .A1 (nx3167), .S0 (nx3248)) ;
    xnor2 ix3847 (.Y (nx3846), .A0 (nx3842), .A1 (nx3185)) ;
    xnor2 ix3843 (.Y (nx3842), .A0 (nx2671), .A1 (nx3840)) ;
    nand02_2x ix3186 (.Y (nx3185), .A0 (input_b[13]), .A1 (input_a[10])) ;
    nand02_2x ix3188 (.Y (nx3187), .A0 (input_b[12]), .A1 (input_a[12])) ;
    xnor2 ix3190 (.Y (nx3189), .A0 (nx3191), .A1 (nx3187)) ;
    xnor2 ix3192 (.Y (nx3191), .A0 (nx3193), .A1 (nx3195)) ;
    mux21_ni ix3194 (.Y (nx3193), .A0 (nx3185), .A1 (nx3179), .S0 (nx3846)) ;
    xnor2 ix3196 (.Y (nx3195), .A0 (nx3197), .A1 (nx3199)) ;
    xnor2 ix3198 (.Y (nx3197), .A0 (nx2667), .A1 (nx2803)) ;
    nand02_2x ix3200 (.Y (nx3199), .A0 (input_b[13]), .A1 (input_a[11])) ;
    xnor2 ix6663 (.Y (nx6662), .A0 (nx6660), .A1 (nx3017)) ;
    xnor2 ix6661 (.Y (nx6660), .A0 (nx3205), .A1 (nx6476)) ;
    mux21_ni ix3206 (.Y (nx3205), .A0 (nx3193), .A1 (nx3199), .S0 (nx3195)) ;
    xnor2 ix6477 (.Y (nx6476), .A0 (nx6474), .A1 (nx3211)) ;
    xnor2 ix6475 (.Y (nx6474), .A0 (nx2665), .A1 (nx6276)) ;
    nand02_2x ix3212 (.Y (nx3211), .A0 (input_b[13]), .A1 (input_a[12])) ;
    nand02_2x ix3214 (.Y (nx3213), .A0 (input_b[12]), .A1 (input_a[14])) ;
    xnor2 ix3216 (.Y (nx3215), .A0 (nx3217), .A1 (nx3213)) ;
    xnor2 ix3218 (.Y (nx3217), .A0 (nx3219), .A1 (nx3221)) ;
    mux21_ni ix3220 (.Y (nx3219), .A0 (nx3211), .A1 (nx3205), .S0 (nx6476)) ;
    xnor2 ix3222 (.Y (nx3221), .A0 (nx3223), .A1 (nx3225)) ;
    xnor2 ix3224 (.Y (nx3223), .A0 (nx2661), .A1 (nx2829)) ;
    nand02_2x ix3226 (.Y (nx3225), .A0 (input_b[13]), .A1 (input_a[13])) ;
    xnor2 ix6643 (.Y (nx6642), .A0 (nx6640), .A1 (nx3011)) ;
    xnor2 ix6641 (.Y (nx6640), .A0 (nx3231), .A1 (nx6456)) ;
    mux21_ni ix3232 (.Y (nx3231), .A0 (nx3219), .A1 (nx3225), .S0 (nx3221)) ;
    xnor2 ix6457 (.Y (nx6456), .A0 (nx6454), .A1 (nx3237)) ;
    xnor2 ix6455 (.Y (nx6454), .A0 (nx2659), .A1 (nx6256)) ;
    nand02_2x ix3238 (.Y (nx3237), .A0 (input_b[13]), .A1 (input_a[14])) ;
    nand02_2x ix3240 (.Y (nx3239), .A0 (input_b[12]), .A1 (input_a[16])) ;
    xnor2 ix3242 (.Y (nx3241), .A0 (nx3243), .A1 (nx3239)) ;
    xnor2 ix3244 (.Y (nx3243), .A0 (nx3245), .A1 (nx3247)) ;
    mux21_ni ix3246 (.Y (nx3245), .A0 (nx3237), .A1 (nx3231), .S0 (nx6456)) ;
    xnor2 ix3248 (.Y (nx3247), .A0 (nx3249), .A1 (nx3251)) ;
    xnor2 ix3250 (.Y (nx3249), .A0 (nx2655), .A1 (nx2855)) ;
    nand02_2x ix3252 (.Y (nx3251), .A0 (input_b[13]), .A1 (input_a[15])) ;
    xnor2 ix6623 (.Y (nx6622), .A0 (nx6620), .A1 (nx3005)) ;
    xnor2 ix6621 (.Y (nx6620), .A0 (nx3257), .A1 (nx6436)) ;
    mux21_ni ix3258 (.Y (nx3257), .A0 (nx3245), .A1 (nx3251), .S0 (nx3247)) ;
    xnor2 ix6437 (.Y (nx6436), .A0 (nx6434), .A1 (nx3263)) ;
    xnor2 ix6435 (.Y (nx6434), .A0 (nx2653), .A1 (nx6236)) ;
    nand02_2x ix3264 (.Y (nx3263), .A0 (input_b[13]), .A1 (input_a[16])) ;
    nand02_2x ix3266 (.Y (nx3265), .A0 (input_b[12]), .A1 (input_a[18])) ;
    xnor2 ix3268 (.Y (nx3267), .A0 (nx3269), .A1 (nx3265)) ;
    xnor2 ix3270 (.Y (nx3269), .A0 (nx3271), .A1 (nx3273)) ;
    mux21_ni ix3272 (.Y (nx3271), .A0 (nx3263), .A1 (nx3257), .S0 (nx6436)) ;
    xnor2 ix3274 (.Y (nx3273), .A0 (nx3275), .A1 (nx3277)) ;
    xnor2 ix3276 (.Y (nx3275), .A0 (nx2649), .A1 (nx2881)) ;
    nand02_2x ix3278 (.Y (nx3277), .A0 (input_b[13]), .A1 (input_a[17])) ;
    xnor2 ix6603 (.Y (nx6602), .A0 (nx6600), .A1 (nx2999)) ;
    xnor2 ix6601 (.Y (nx6600), .A0 (nx3283), .A1 (nx6416)) ;
    mux21_ni ix3284 (.Y (nx3283), .A0 (nx3271), .A1 (nx3277), .S0 (nx3273)) ;
    xnor2 ix6417 (.Y (nx6416), .A0 (nx6414), .A1 (nx3289)) ;
    xnor2 ix6415 (.Y (nx6414), .A0 (nx2647), .A1 (nx6216)) ;
    nand02_2x ix3290 (.Y (nx3289), .A0 (input_b[13]), .A1 (input_a[18])) ;
    nand02_2x ix3292 (.Y (nx3291), .A0 (input_b[12]), .A1 (input_a[20])) ;
    xnor2 ix3294 (.Y (nx3293), .A0 (nx3295), .A1 (nx3291)) ;
    xnor2 ix3296 (.Y (nx3295), .A0 (nx3297), .A1 (nx3299)) ;
    mux21_ni ix3298 (.Y (nx3297), .A0 (nx3289), .A1 (nx3283), .S0 (nx6416)) ;
    xnor2 ix3300 (.Y (nx3299), .A0 (nx3301), .A1 (nx3303)) ;
    xnor2 ix3302 (.Y (nx3301), .A0 (nx2643), .A1 (nx2907)) ;
    nand02_2x ix3304 (.Y (nx3303), .A0 (input_b[13]), .A1 (input_a[19])) ;
    xnor2 ix6583 (.Y (nx6582), .A0 (nx6580), .A1 (nx2993)) ;
    xnor2 ix6581 (.Y (nx6580), .A0 (nx3309), .A1 (nx6396)) ;
    mux21_ni ix3310 (.Y (nx3309), .A0 (nx3297), .A1 (nx3303), .S0 (nx3299)) ;
    xnor2 ix6397 (.Y (nx6396), .A0 (nx6394), .A1 (nx3315)) ;
    xnor2 ix6395 (.Y (nx6394), .A0 (nx2641), .A1 (nx6196)) ;
    nand02_2x ix3316 (.Y (nx3315), .A0 (input_b[13]), .A1 (input_a[20])) ;
    nand02_2x ix3318 (.Y (nx3317), .A0 (input_b[12]), .A1 (input_a[22])) ;
    xnor2 ix3320 (.Y (nx3319), .A0 (nx3321), .A1 (nx3317)) ;
    xnor2 ix3322 (.Y (nx3321), .A0 (nx3323), .A1 (nx3325)) ;
    mux21_ni ix3324 (.Y (nx3323), .A0 (nx3315), .A1 (nx3309), .S0 (nx6396)) ;
    xnor2 ix3326 (.Y (nx3325), .A0 (nx3327), .A1 (nx3329)) ;
    xnor2 ix3328 (.Y (nx3327), .A0 (nx2637), .A1 (nx2933)) ;
    nand02_2x ix3330 (.Y (nx3329), .A0 (input_b[13]), .A1 (input_a[21])) ;
    xnor2 ix3332 (.Y (nx3331), .A0 (input_b[12]), .A1 (nx6560)) ;
    xnor2 ix6561 (.Y (nx6560), .A0 (nx3335), .A1 (nx6376)) ;
    mux21_ni ix3336 (.Y (nx3335), .A0 (nx3323), .A1 (nx3329), .S0 (nx3325)) ;
    xnor2 ix6377 (.Y (nx6376), .A0 (nx6374), .A1 (nx3341)) ;
    xnor2 ix6375 (.Y (nx6374), .A0 (nx2635), .A1 (nx6176)) ;
    nand02_2x ix3342 (.Y (nx3341), .A0 (input_b[13]), .A1 (input_a[22])) ;
    mux21_ni ix7865 (.Y (nx7864), .A0 (nx7062), .A1 (nx7860), .S0 (nx7196)) ;
    mux21_ni ix3350 (.Y (nx3349), .A0 (nx3351), .A1 (nx3677), .S0 (nx3679)) ;
    mux21_ni ix3352 (.Y (nx3351), .A0 (nx3353), .A1 (nx3355), .S0 (nx6932)) ;
    nand02_2x ix3354 (.Y (nx3353), .A0 (input_b[10]), .A1 (input_a[21])) ;
    mux21_ni ix3356 (.Y (nx3355), .A0 (nx3357), .A1 (nx3651), .S0 (nx3653)) ;
    mux21_ni ix3358 (.Y (nx3357), .A0 (nx3359), .A1 (nx3361), .S0 (nx6952)) ;
    nand02_2x ix3360 (.Y (nx3359), .A0 (input_b[10]), .A1 (input_a[19])) ;
    mux21_ni ix3362 (.Y (nx3361), .A0 (nx3363), .A1 (nx3625), .S0 (nx3627)) ;
    mux21_ni ix3364 (.Y (nx3363), .A0 (nx3365), .A1 (nx3367), .S0 (nx6972)) ;
    nand02_2x ix3366 (.Y (nx3365), .A0 (input_b[10]), .A1 (input_a[17])) ;
    mux21_ni ix3368 (.Y (nx3367), .A0 (nx3369), .A1 (nx3599), .S0 (nx3601)) ;
    mux21_ni ix3370 (.Y (nx3369), .A0 (nx3371), .A1 (nx3373), .S0 (nx6992)) ;
    nand02_2x ix3372 (.Y (nx3371), .A0 (input_b[10]), .A1 (input_a[15])) ;
    mux21_ni ix3374 (.Y (nx3373), .A0 (nx3375), .A1 (nx3573), .S0 (nx3575)) ;
    mux21_ni ix3376 (.Y (nx3375), .A0 (nx3377), .A1 (nx3379), .S0 (nx3864)) ;
    nand02_2x ix3378 (.Y (nx3377), .A0 (input_b[10]), .A1 (input_a[13])) ;
    mux21_ni ix3380 (.Y (nx3379), .A0 (nx3381), .A1 (nx3383), .S0 (nx3266)) ;
    nand02_2x ix3382 (.Y (nx3381), .A0 (input_b[10]), .A1 (input_a[12])) ;
    mux21_ni ix3384 (.Y (nx3383), .A0 (nx3385), .A1 (nx3535), .S0 (nx3537)) ;
    mux21_ni ix3386 (.Y (nx3385), .A0 (nx3387), .A1 (nx3521), .S0 (nx3523)) ;
    mux21_ni ix3388 (.Y (nx3387), .A0 (nx3389), .A1 (nx3507), .S0 (nx3509)) ;
    mux21_ni ix3390 (.Y (nx3389), .A0 (nx3391), .A1 (nx3493), .S0 (nx3495)) ;
    mux21_ni ix3392 (.Y (nx3391), .A0 (nx3393), .A1 (nx3479), .S0 (nx3481)) ;
    mux21_ni ix3394 (.Y (nx3393), .A0 (nx3395), .A1 (nx3465), .S0 (nx3467)) ;
    mux21_ni ix3396 (.Y (nx3395), .A0 (nx3397), .A1 (nx3451), .S0 (nx3453)) ;
    mux21_ni ix3398 (.Y (nx3397), .A0 (nx3399), .A1 (nx3435), .S0 (nx3437)) ;
    mux21_ni ix3400 (.Y (nx3399), .A0 (nx3401), .A1 (nx3419), .S0 (nx3421)) ;
    mux21_ni ix3402 (.Y (nx3401), .A0 (nx3403), .A1 (nx3405), .S0 (nx292)) ;
    nand02_2x ix3404 (.Y (nx3403), .A0 (input_b[10]), .A1 (input_a[2])) ;
    xnor2 ix293 (.Y (nx292), .A0 (nx290), .A1 (nx3403)) ;
    inv02 ix3414 (.Y (nx3413), .A (input_b[11])) ;
    inv02 ix3416 (.Y (nx3415), .A (input_b[12])) ;
    aoi22 ix3418 (.Y (nx3417), .A0 (input_b[12]), .A1 (input_a[0]), .B0 (
          input_b[11]), .B1 (input_a[1])) ;
    nand02_2x ix3420 (.Y (nx3419), .A0 (input_b[10]), .A1 (input_a[3])) ;
    xnor2 ix3422 (.Y (nx3421), .A0 (nx3423), .A1 (nx3419)) ;
    xnor2 ix327 (.Y (nx326), .A0 (nx322), .A1 (nx3433)) ;
    aoi22 ix3432 (.Y (nx3431), .A0 (input_b[13]), .A1 (input_a[0]), .B0 (
          input_b[12]), .B1 (input_a[1])) ;
    nand02_2x ix3434 (.Y (nx3433), .A0 (input_b[11]), .A1 (input_a[2])) ;
    nand02_2x ix3436 (.Y (nx3435), .A0 (input_b[10]), .A1 (input_a[4])) ;
    xnor2 ix3438 (.Y (nx3437), .A0 (nx3439), .A1 (nx3435)) ;
    xnor2 ix3440 (.Y (nx3439), .A0 (nx3441), .A1 (nx3445)) ;
    mux21_ni ix3442 (.Y (nx3441), .A0 (nx3433), .A1 (nx3443), .S0 (nx326)) ;
    xnor2 ix3446 (.Y (nx3445), .A0 (nx3447), .A1 (nx3449)) ;
    nand02_2x ix3450 (.Y (nx3449), .A0 (input_b[11]), .A1 (input_a[3])) ;
    nand02_2x ix3452 (.Y (nx3451), .A0 (input_b[10]), .A1 (input_a[5])) ;
    xnor2 ix3454 (.Y (nx3453), .A0 (nx3455), .A1 (nx3451)) ;
    xnor2 ix3456 (.Y (nx3455), .A0 (nx3457), .A1 (nx3459)) ;
    mux21_ni ix3458 (.Y (nx3457), .A0 (nx3441), .A1 (nx3449), .S0 (nx3445)) ;
    xnor2 ix3460 (.Y (nx3459), .A0 (nx3461), .A1 (nx3463)) ;
    xnor2 ix3462 (.Y (nx3461), .A0 (nx3043), .A1 (nx3063)) ;
    nand02_2x ix3464 (.Y (nx3463), .A0 (input_b[11]), .A1 (input_a[4])) ;
    nand02_2x ix3466 (.Y (nx3465), .A0 (input_b[10]), .A1 (input_a[6])) ;
    xnor2 ix3468 (.Y (nx3467), .A0 (nx3469), .A1 (nx3465)) ;
    xnor2 ix3470 (.Y (nx3469), .A0 (nx3471), .A1 (nx3473)) ;
    mux21_ni ix3472 (.Y (nx3471), .A0 (nx3457), .A1 (nx3463), .S0 (nx3459)) ;
    xnor2 ix3474 (.Y (nx3473), .A0 (nx3475), .A1 (nx3477)) ;
    xnor2 ix3476 (.Y (nx3475), .A0 (nx3041), .A1 (nx3079)) ;
    nand02_2x ix3478 (.Y (nx3477), .A0 (input_b[11]), .A1 (input_a[5])) ;
    nand02_2x ix3480 (.Y (nx3479), .A0 (input_b[10]), .A1 (input_a[7])) ;
    xnor2 ix3482 (.Y (nx3481), .A0 (nx3483), .A1 (nx3479)) ;
    xnor2 ix3484 (.Y (nx3483), .A0 (nx3485), .A1 (nx3487)) ;
    mux21_ni ix3486 (.Y (nx3485), .A0 (nx3471), .A1 (nx3477), .S0 (nx3473)) ;
    xnor2 ix3488 (.Y (nx3487), .A0 (nx3489), .A1 (nx3491)) ;
    xnor2 ix3490 (.Y (nx3489), .A0 (nx3039), .A1 (nx3095)) ;
    nand02_2x ix3492 (.Y (nx3491), .A0 (input_b[11]), .A1 (input_a[6])) ;
    nand02_2x ix3494 (.Y (nx3493), .A0 (input_b[10]), .A1 (input_a[8])) ;
    xnor2 ix3496 (.Y (nx3495), .A0 (nx3497), .A1 (nx3493)) ;
    xnor2 ix3498 (.Y (nx3497), .A0 (nx3499), .A1 (nx3501)) ;
    mux21_ni ix3500 (.Y (nx3499), .A0 (nx3485), .A1 (nx3491), .S0 (nx3487)) ;
    xnor2 ix3502 (.Y (nx3501), .A0 (nx3503), .A1 (nx3505)) ;
    xnor2 ix3504 (.Y (nx3503), .A0 (nx3037), .A1 (nx3109)) ;
    nand02_2x ix3506 (.Y (nx3505), .A0 (input_b[11]), .A1 (input_a[7])) ;
    nand02_2x ix3508 (.Y (nx3507), .A0 (input_b[10]), .A1 (input_a[9])) ;
    xnor2 ix3510 (.Y (nx3509), .A0 (nx3511), .A1 (nx3507)) ;
    xnor2 ix3512 (.Y (nx3511), .A0 (nx3513), .A1 (nx3515)) ;
    mux21_ni ix3514 (.Y (nx3513), .A0 (nx3499), .A1 (nx3505), .S0 (nx3501)) ;
    xnor2 ix3516 (.Y (nx3515), .A0 (nx3517), .A1 (nx3519)) ;
    xnor2 ix3518 (.Y (nx3517), .A0 (nx3035), .A1 (nx3123)) ;
    nand02_2x ix3520 (.Y (nx3519), .A0 (input_b[11]), .A1 (input_a[8])) ;
    nand02_2x ix3522 (.Y (nx3521), .A0 (input_b[10]), .A1 (input_a[10])) ;
    xnor2 ix3524 (.Y (nx3523), .A0 (nx3525), .A1 (nx3521)) ;
    xnor2 ix3526 (.Y (nx3525), .A0 (nx3527), .A1 (nx3529)) ;
    mux21_ni ix3528 (.Y (nx3527), .A0 (nx3513), .A1 (nx3519), .S0 (nx3515)) ;
    xnor2 ix3530 (.Y (nx3529), .A0 (nx3531), .A1 (nx3533)) ;
    xnor2 ix3532 (.Y (nx3531), .A0 (nx3033), .A1 (nx3137)) ;
    nand02_2x ix3534 (.Y (nx3533), .A0 (input_b[11]), .A1 (input_a[9])) ;
    nand02_2x ix3536 (.Y (nx3535), .A0 (input_b[10]), .A1 (input_a[11])) ;
    xnor2 ix3538 (.Y (nx3537), .A0 (nx3539), .A1 (nx3535)) ;
    xnor2 ix3540 (.Y (nx3539), .A0 (nx3541), .A1 (nx3543)) ;
    mux21_ni ix3542 (.Y (nx3541), .A0 (nx3527), .A1 (nx3533), .S0 (nx3529)) ;
    xnor2 ix3544 (.Y (nx3543), .A0 (nx3545), .A1 (nx3547)) ;
    xnor2 ix3546 (.Y (nx3545), .A0 (nx3031), .A1 (nx3151)) ;
    nand02_2x ix3548 (.Y (nx3547), .A0 (input_b[11]), .A1 (input_a[10])) ;
    xnor2 ix3267 (.Y (nx3266), .A0 (nx3262), .A1 (nx3381)) ;
    xnor2 ix3263 (.Y (nx3262), .A0 (nx3553), .A1 (nx3260)) ;
    mux21_ni ix3554 (.Y (nx3553), .A0 (nx3541), .A1 (nx3547), .S0 (nx3543)) ;
    xnor2 ix3261 (.Y (nx3260), .A0 (nx3256), .A1 (nx3559)) ;
    xnor2 ix3257 (.Y (nx3256), .A0 (nx3029), .A1 (nx3254)) ;
    nand02_2x ix3560 (.Y (nx3559), .A0 (input_b[11]), .A1 (input_a[11])) ;
    xnor2 ix3865 (.Y (nx3864), .A0 (nx3860), .A1 (nx3377)) ;
    xnor2 ix3861 (.Y (nx3860), .A0 (nx3565), .A1 (nx3858)) ;
    mux21_ni ix3566 (.Y (nx3565), .A0 (nx3559), .A1 (nx3553), .S0 (nx3260)) ;
    xnor2 ix3859 (.Y (nx3858), .A0 (nx3854), .A1 (nx3571)) ;
    xnor2 ix3855 (.Y (nx3854), .A0 (nx3025), .A1 (nx3852)) ;
    nand02_2x ix3572 (.Y (nx3571), .A0 (input_b[11]), .A1 (input_a[12])) ;
    nand02_2x ix3574 (.Y (nx3573), .A0 (input_b[10]), .A1 (input_a[14])) ;
    xnor2 ix3576 (.Y (nx3575), .A0 (nx3577), .A1 (nx3573)) ;
    xnor2 ix3578 (.Y (nx3577), .A0 (nx3579), .A1 (nx3581)) ;
    mux21_ni ix3580 (.Y (nx3579), .A0 (nx3571), .A1 (nx3565), .S0 (nx3858)) ;
    xnor2 ix3582 (.Y (nx3581), .A0 (nx3583), .A1 (nx3585)) ;
    xnor2 ix3584 (.Y (nx3583), .A0 (nx3021), .A1 (nx3189)) ;
    nand02_2x ix3586 (.Y (nx3585), .A0 (input_b[11]), .A1 (input_a[13])) ;
    xnor2 ix6993 (.Y (nx6992), .A0 (nx6990), .A1 (nx3371)) ;
    xnor2 ix6991 (.Y (nx6990), .A0 (nx3591), .A1 (nx6834)) ;
    mux21_ni ix3592 (.Y (nx3591), .A0 (nx3579), .A1 (nx3585), .S0 (nx3581)) ;
    xnor2 ix6835 (.Y (nx6834), .A0 (nx6832), .A1 (nx3597)) ;
    xnor2 ix6833 (.Y (nx6832), .A0 (nx3019), .A1 (nx6662)) ;
    nand02_2x ix3598 (.Y (nx3597), .A0 (input_b[11]), .A1 (input_a[14])) ;
    nand02_2x ix3600 (.Y (nx3599), .A0 (input_b[10]), .A1 (input_a[16])) ;
    xnor2 ix3602 (.Y (nx3601), .A0 (nx3603), .A1 (nx3599)) ;
    xnor2 ix3604 (.Y (nx3603), .A0 (nx3605), .A1 (nx3607)) ;
    mux21_ni ix3606 (.Y (nx3605), .A0 (nx3597), .A1 (nx3591), .S0 (nx6834)) ;
    xnor2 ix3608 (.Y (nx3607), .A0 (nx3609), .A1 (nx3611)) ;
    xnor2 ix3610 (.Y (nx3609), .A0 (nx3015), .A1 (nx3215)) ;
    nand02_2x ix3612 (.Y (nx3611), .A0 (input_b[11]), .A1 (input_a[15])) ;
    xnor2 ix6973 (.Y (nx6972), .A0 (nx6970), .A1 (nx3365)) ;
    xnor2 ix6971 (.Y (nx6970), .A0 (nx3617), .A1 (nx6814)) ;
    mux21_ni ix3618 (.Y (nx3617), .A0 (nx3605), .A1 (nx3611), .S0 (nx3607)) ;
    xnor2 ix6815 (.Y (nx6814), .A0 (nx6812), .A1 (nx3623)) ;
    xnor2 ix6813 (.Y (nx6812), .A0 (nx3013), .A1 (nx6642)) ;
    nand02_2x ix3624 (.Y (nx3623), .A0 (input_b[11]), .A1 (input_a[16])) ;
    nand02_2x ix3626 (.Y (nx3625), .A0 (input_b[10]), .A1 (input_a[18])) ;
    xnor2 ix3628 (.Y (nx3627), .A0 (nx3629), .A1 (nx3625)) ;
    xnor2 ix3630 (.Y (nx3629), .A0 (nx3631), .A1 (nx3633)) ;
    mux21_ni ix3632 (.Y (nx3631), .A0 (nx3623), .A1 (nx3617), .S0 (nx6814)) ;
    xnor2 ix3634 (.Y (nx3633), .A0 (nx3635), .A1 (nx3637)) ;
    xnor2 ix3636 (.Y (nx3635), .A0 (nx3009), .A1 (nx3241)) ;
    nand02_2x ix3638 (.Y (nx3637), .A0 (input_b[11]), .A1 (input_a[17])) ;
    xnor2 ix6953 (.Y (nx6952), .A0 (nx6950), .A1 (nx3359)) ;
    xnor2 ix6951 (.Y (nx6950), .A0 (nx3643), .A1 (nx6794)) ;
    mux21_ni ix3644 (.Y (nx3643), .A0 (nx3631), .A1 (nx3637), .S0 (nx3633)) ;
    xnor2 ix6795 (.Y (nx6794), .A0 (nx6792), .A1 (nx3649)) ;
    xnor2 ix6793 (.Y (nx6792), .A0 (nx3007), .A1 (nx6622)) ;
    nand02_2x ix3650 (.Y (nx3649), .A0 (input_b[11]), .A1 (input_a[18])) ;
    nand02_2x ix3652 (.Y (nx3651), .A0 (input_b[10]), .A1 (input_a[20])) ;
    xnor2 ix3654 (.Y (nx3653), .A0 (nx3655), .A1 (nx3651)) ;
    xnor2 ix3656 (.Y (nx3655), .A0 (nx3657), .A1 (nx3659)) ;
    mux21_ni ix3658 (.Y (nx3657), .A0 (nx3649), .A1 (nx3643), .S0 (nx6794)) ;
    xnor2 ix3660 (.Y (nx3659), .A0 (nx3661), .A1 (nx3663)) ;
    xnor2 ix3662 (.Y (nx3661), .A0 (nx3003), .A1 (nx3267)) ;
    nand02_2x ix3664 (.Y (nx3663), .A0 (input_b[11]), .A1 (input_a[19])) ;
    xnor2 ix6933 (.Y (nx6932), .A0 (nx6930), .A1 (nx3353)) ;
    xnor2 ix6931 (.Y (nx6930), .A0 (nx3669), .A1 (nx6774)) ;
    mux21_ni ix3670 (.Y (nx3669), .A0 (nx3657), .A1 (nx3663), .S0 (nx3659)) ;
    xnor2 ix6775 (.Y (nx6774), .A0 (nx6772), .A1 (nx3675)) ;
    xnor2 ix6773 (.Y (nx6772), .A0 (nx3001), .A1 (nx6602)) ;
    nand02_2x ix3676 (.Y (nx3675), .A0 (input_b[11]), .A1 (input_a[20])) ;
    nand02_2x ix3678 (.Y (nx3677), .A0 (input_b[10]), .A1 (input_a[22])) ;
    xnor2 ix3680 (.Y (nx3679), .A0 (nx3681), .A1 (nx3677)) ;
    xnor2 ix3682 (.Y (nx3681), .A0 (nx3683), .A1 (nx3685)) ;
    mux21_ni ix3684 (.Y (nx3683), .A0 (nx3675), .A1 (nx3669), .S0 (nx6774)) ;
    xnor2 ix3686 (.Y (nx3685), .A0 (nx3687), .A1 (nx3689)) ;
    xnor2 ix3688 (.Y (nx3687), .A0 (nx2997), .A1 (nx3293)) ;
    nand02_2x ix3690 (.Y (nx3689), .A0 (input_b[11]), .A1 (input_a[21])) ;
    xnor2 ix3692 (.Y (nx3691), .A0 (input_b[10]), .A1 (nx6910)) ;
    xnor2 ix6911 (.Y (nx6910), .A0 (nx3695), .A1 (nx6754)) ;
    mux21_ni ix3696 (.Y (nx3695), .A0 (nx3683), .A1 (nx3689), .S0 (nx3685)) ;
    xnor2 ix6755 (.Y (nx6754), .A0 (nx6752), .A1 (nx3701)) ;
    xnor2 ix6753 (.Y (nx6752), .A0 (nx2995), .A1 (nx6582)) ;
    nand02_2x ix3702 (.Y (nx3701), .A0 (input_b[11]), .A1 (input_a[22])) ;
    mux21_ni ix7861 (.Y (nx7860), .A0 (nx7856), .A1 (nx7202), .S0 (nx5591)) ;
    xnor2 ix3708 (.Y (nx3707), .A0 (nx3709), .A1 (nx4051)) ;
    mux21_ni ix3710 (.Y (nx3709), .A0 (nx3711), .A1 (nx4037), .S0 (nx4039)) ;
    mux21_ni ix3712 (.Y (nx3711), .A0 (nx3713), .A1 (nx3715), .S0 (nx7226)) ;
    nand02_2x ix3714 (.Y (nx3713), .A0 (input_b[8]), .A1 (input_a[21])) ;
    mux21_ni ix3716 (.Y (nx3715), .A0 (nx3717), .A1 (nx4011), .S0 (nx4013)) ;
    mux21_ni ix3718 (.Y (nx3717), .A0 (nx3719), .A1 (nx3721), .S0 (nx7246)) ;
    nand02_2x ix3720 (.Y (nx3719), .A0 (input_b[8]), .A1 (input_a[19])) ;
    mux21_ni ix3722 (.Y (nx3721), .A0 (nx3723), .A1 (nx3985), .S0 (nx3987)) ;
    mux21_ni ix3724 (.Y (nx3723), .A0 (nx3725), .A1 (nx3727), .S0 (nx7266)) ;
    nand02_2x ix3726 (.Y (nx3725), .A0 (input_b[8]), .A1 (input_a[17])) ;
    mux21_ni ix3728 (.Y (nx3727), .A0 (nx3729), .A1 (nx3959), .S0 (nx3961)) ;
    mux21_ni ix3730 (.Y (nx3729), .A0 (nx3731), .A1 (nx3733), .S0 (nx3876)) ;
    nand02_2x ix3732 (.Y (nx3731), .A0 (input_b[8]), .A1 (input_a[15])) ;
    mux21_ni ix3734 (.Y (nx3733), .A0 (nx3735), .A1 (nx3737), .S0 (nx3278)) ;
    nand02_2x ix3736 (.Y (nx3735), .A0 (input_b[8]), .A1 (input_a[14])) ;
    mux21_ni ix3738 (.Y (nx3737), .A0 (nx3739), .A1 (nx3921), .S0 (nx3923)) ;
    mux21_ni ix3740 (.Y (nx3739), .A0 (nx3741), .A1 (nx3907), .S0 (nx3909)) ;
    mux21_ni ix3742 (.Y (nx3741), .A0 (nx3743), .A1 (nx3893), .S0 (nx3895)) ;
    mux21_ni ix3744 (.Y (nx3743), .A0 (nx3745), .A1 (nx3879), .S0 (nx3881)) ;
    mux21_ni ix3746 (.Y (nx3745), .A0 (nx3747), .A1 (nx3865), .S0 (nx3867)) ;
    mux21_ni ix3748 (.Y (nx3747), .A0 (nx3749), .A1 (nx3851), .S0 (nx3853)) ;
    mux21_ni ix3750 (.Y (nx3749), .A0 (nx3751), .A1 (nx3837), .S0 (nx3839)) ;
    mux21_ni ix3752 (.Y (nx3751), .A0 (nx3753), .A1 (nx3823), .S0 (nx3825)) ;
    mux21_ni ix3754 (.Y (nx3753), .A0 (nx3755), .A1 (nx3809), .S0 (nx3811)) ;
    mux21_ni ix3756 (.Y (nx3755), .A0 (nx3757), .A1 (nx3793), .S0 (nx3795)) ;
    mux21_ni ix3758 (.Y (nx3757), .A0 (nx3759), .A1 (nx3777), .S0 (nx3779)) ;
    mux21_ni ix3760 (.Y (nx3759), .A0 (nx3761), .A1 (nx3763), .S0 (nx492)) ;
    nand02_2x ix3762 (.Y (nx3761), .A0 (input_b[8]), .A1 (input_a[2])) ;
    xnor2 ix493 (.Y (nx492), .A0 (nx490), .A1 (nx3761)) ;
    inv02 ix3772 (.Y (nx3771), .A (input_b[9])) ;
    inv02 ix3774 (.Y (nx3773), .A (input_b[10])) ;
    aoi22 ix3776 (.Y (nx3775), .A0 (input_b[10]), .A1 (input_a[0]), .B0 (
          input_b[9]), .B1 (input_a[1])) ;
    nand02_2x ix3778 (.Y (nx3777), .A0 (input_b[8]), .A1 (input_a[3])) ;
    xnor2 ix3780 (.Y (nx3779), .A0 (nx3781), .A1 (nx3777)) ;
    xnor2 ix365 (.Y (nx364), .A0 (nx362), .A1 (nx3791)) ;
    aoi22 ix3790 (.Y (nx3789), .A0 (input_b[11]), .A1 (input_a[0]), .B0 (
          input_b[10]), .B1 (input_a[1])) ;
    nand02_2x ix3792 (.Y (nx3791), .A0 (input_b[9]), .A1 (input_a[2])) ;
    nand02_2x ix3794 (.Y (nx3793), .A0 (input_b[8]), .A1 (input_a[4])) ;
    xnor2 ix3796 (.Y (nx3795), .A0 (nx3797), .A1 (nx3793)) ;
    xnor2 ix3798 (.Y (nx3797), .A0 (nx3799), .A1 (nx3803)) ;
    mux21_ni ix3800 (.Y (nx3799), .A0 (nx3791), .A1 (nx3801), .S0 (nx364)) ;
    xnor2 ix3804 (.Y (nx3803), .A0 (nx3805), .A1 (nx3807)) ;
    nand02_2x ix3808 (.Y (nx3807), .A0 (input_b[9]), .A1 (input_a[3])) ;
    nand02_2x ix3810 (.Y (nx3809), .A0 (input_b[8]), .A1 (input_a[5])) ;
    xnor2 ix3812 (.Y (nx3811), .A0 (nx3813), .A1 (nx3809)) ;
    xnor2 ix3814 (.Y (nx3813), .A0 (nx3815), .A1 (nx3817)) ;
    mux21_ni ix3816 (.Y (nx3815), .A0 (nx3799), .A1 (nx3807), .S0 (nx3803)) ;
    xnor2 ix3818 (.Y (nx3817), .A0 (nx3819), .A1 (nx3821)) ;
    xnor2 ix3820 (.Y (nx3819), .A0 (nx3401), .A1 (nx3421)) ;
    nand02_2x ix3822 (.Y (nx3821), .A0 (input_b[9]), .A1 (input_a[4])) ;
    nand02_2x ix3824 (.Y (nx3823), .A0 (input_b[8]), .A1 (input_a[6])) ;
    xnor2 ix3826 (.Y (nx3825), .A0 (nx3827), .A1 (nx3823)) ;
    xnor2 ix3828 (.Y (nx3827), .A0 (nx3829), .A1 (nx3831)) ;
    mux21_ni ix3830 (.Y (nx3829), .A0 (nx3815), .A1 (nx3821), .S0 (nx3817)) ;
    xnor2 ix3832 (.Y (nx3831), .A0 (nx3833), .A1 (nx3835)) ;
    xnor2 ix3834 (.Y (nx3833), .A0 (nx3399), .A1 (nx3437)) ;
    nand02_2x ix3836 (.Y (nx3835), .A0 (input_b[9]), .A1 (input_a[5])) ;
    nand02_2x ix3838 (.Y (nx3837), .A0 (input_b[8]), .A1 (input_a[7])) ;
    xnor2 ix3840 (.Y (nx3839), .A0 (nx3841), .A1 (nx3837)) ;
    xnor2 ix3842 (.Y (nx3841), .A0 (nx3843), .A1 (nx3845)) ;
    mux21_ni ix3844 (.Y (nx3843), .A0 (nx3829), .A1 (nx3835), .S0 (nx3831)) ;
    xnor2 ix3846 (.Y (nx3845), .A0 (nx3847), .A1 (nx3849)) ;
    xnor2 ix3848 (.Y (nx3847), .A0 (nx3397), .A1 (nx3453)) ;
    nand02_2x ix3850 (.Y (nx3849), .A0 (input_b[9]), .A1 (input_a[6])) ;
    nand02_2x ix3852 (.Y (nx3851), .A0 (input_b[8]), .A1 (input_a[8])) ;
    xnor2 ix3854 (.Y (nx3853), .A0 (nx3855), .A1 (nx3851)) ;
    xnor2 ix3856 (.Y (nx3855), .A0 (nx3857), .A1 (nx3859)) ;
    mux21_ni ix3858 (.Y (nx3857), .A0 (nx3843), .A1 (nx3849), .S0 (nx3845)) ;
    xnor2 ix3860 (.Y (nx3859), .A0 (nx3861), .A1 (nx3863)) ;
    xnor2 ix3862 (.Y (nx3861), .A0 (nx3395), .A1 (nx3467)) ;
    nand02_2x ix3864 (.Y (nx3863), .A0 (input_b[9]), .A1 (input_a[7])) ;
    nand02_2x ix3866 (.Y (nx3865), .A0 (input_b[8]), .A1 (input_a[9])) ;
    xnor2 ix3868 (.Y (nx3867), .A0 (nx3869), .A1 (nx3865)) ;
    xnor2 ix3870 (.Y (nx3869), .A0 (nx3871), .A1 (nx3873)) ;
    mux21_ni ix3872 (.Y (nx3871), .A0 (nx3857), .A1 (nx3863), .S0 (nx3859)) ;
    xnor2 ix3874 (.Y (nx3873), .A0 (nx3875), .A1 (nx3877)) ;
    xnor2 ix3876 (.Y (nx3875), .A0 (nx3393), .A1 (nx3481)) ;
    nand02_2x ix3878 (.Y (nx3877), .A0 (input_b[9]), .A1 (input_a[8])) ;
    nand02_2x ix3880 (.Y (nx3879), .A0 (input_b[8]), .A1 (input_a[10])) ;
    xnor2 ix3882 (.Y (nx3881), .A0 (nx3883), .A1 (nx3879)) ;
    xnor2 ix3884 (.Y (nx3883), .A0 (nx3885), .A1 (nx3887)) ;
    mux21_ni ix3886 (.Y (nx3885), .A0 (nx3871), .A1 (nx3877), .S0 (nx3873)) ;
    xnor2 ix3888 (.Y (nx3887), .A0 (nx3889), .A1 (nx3891)) ;
    xnor2 ix3890 (.Y (nx3889), .A0 (nx3391), .A1 (nx3495)) ;
    nand02_2x ix3892 (.Y (nx3891), .A0 (input_b[9]), .A1 (input_a[9])) ;
    nand02_2x ix3894 (.Y (nx3893), .A0 (input_b[8]), .A1 (input_a[11])) ;
    xnor2 ix3896 (.Y (nx3895), .A0 (nx3897), .A1 (nx3893)) ;
    xnor2 ix3898 (.Y (nx3897), .A0 (nx3899), .A1 (nx3901)) ;
    mux21_ni ix3900 (.Y (nx3899), .A0 (nx3885), .A1 (nx3891), .S0 (nx3887)) ;
    xnor2 ix3902 (.Y (nx3901), .A0 (nx3903), .A1 (nx3905)) ;
    xnor2 ix3904 (.Y (nx3903), .A0 (nx3389), .A1 (nx3509)) ;
    nand02_2x ix3906 (.Y (nx3905), .A0 (input_b[9]), .A1 (input_a[10])) ;
    nand02_2x ix3908 (.Y (nx3907), .A0 (input_b[8]), .A1 (input_a[12])) ;
    xnor2 ix3910 (.Y (nx3909), .A0 (nx3911), .A1 (nx3907)) ;
    xnor2 ix3912 (.Y (nx3911), .A0 (nx3913), .A1 (nx3915)) ;
    mux21_ni ix3914 (.Y (nx3913), .A0 (nx3899), .A1 (nx3905), .S0 (nx3901)) ;
    xnor2 ix3916 (.Y (nx3915), .A0 (nx3917), .A1 (nx3919)) ;
    xnor2 ix3918 (.Y (nx3917), .A0 (nx3387), .A1 (nx3523)) ;
    nand02_2x ix3920 (.Y (nx3919), .A0 (input_b[9]), .A1 (input_a[11])) ;
    nand02_2x ix3922 (.Y (nx3921), .A0 (input_b[8]), .A1 (input_a[13])) ;
    xnor2 ix3924 (.Y (nx3923), .A0 (nx3925), .A1 (nx3921)) ;
    xnor2 ix3926 (.Y (nx3925), .A0 (nx3927), .A1 (nx3929)) ;
    mux21_ni ix3928 (.Y (nx3927), .A0 (nx3913), .A1 (nx3919), .S0 (nx3915)) ;
    xnor2 ix3930 (.Y (nx3929), .A0 (nx3931), .A1 (nx3933)) ;
    xnor2 ix3932 (.Y (nx3931), .A0 (nx3385), .A1 (nx3537)) ;
    nand02_2x ix3934 (.Y (nx3933), .A0 (input_b[9]), .A1 (input_a[12])) ;
    xnor2 ix3279 (.Y (nx3278), .A0 (nx3274), .A1 (nx3735)) ;
    xnor2 ix3275 (.Y (nx3274), .A0 (nx3939), .A1 (nx3272)) ;
    mux21_ni ix3940 (.Y (nx3939), .A0 (nx3927), .A1 (nx3933), .S0 (nx3929)) ;
    xnor2 ix3273 (.Y (nx3272), .A0 (nx3268), .A1 (nx3945)) ;
    xnor2 ix3269 (.Y (nx3268), .A0 (nx3383), .A1 (nx3266)) ;
    nand02_2x ix3946 (.Y (nx3945), .A0 (input_b[9]), .A1 (input_a[13])) ;
    xnor2 ix3877 (.Y (nx3876), .A0 (nx3872), .A1 (nx3731)) ;
    xnor2 ix3873 (.Y (nx3872), .A0 (nx3951), .A1 (nx3870)) ;
    mux21_ni ix3952 (.Y (nx3951), .A0 (nx3945), .A1 (nx3939), .S0 (nx3272)) ;
    xnor2 ix3871 (.Y (nx3870), .A0 (nx3866), .A1 (nx3957)) ;
    xnor2 ix3867 (.Y (nx3866), .A0 (nx3379), .A1 (nx3864)) ;
    nand02_2x ix3958 (.Y (nx3957), .A0 (input_b[9]), .A1 (input_a[14])) ;
    nand02_2x ix3960 (.Y (nx3959), .A0 (input_b[8]), .A1 (input_a[16])) ;
    xnor2 ix3962 (.Y (nx3961), .A0 (nx3963), .A1 (nx3959)) ;
    xnor2 ix3964 (.Y (nx3963), .A0 (nx3965), .A1 (nx3967)) ;
    mux21_ni ix3966 (.Y (nx3965), .A0 (nx3957), .A1 (nx3951), .S0 (nx3870)) ;
    xnor2 ix3968 (.Y (nx3967), .A0 (nx3969), .A1 (nx3971)) ;
    xnor2 ix3970 (.Y (nx3969), .A0 (nx3375), .A1 (nx3575)) ;
    nand02_2x ix3972 (.Y (nx3971), .A0 (input_b[9]), .A1 (input_a[15])) ;
    xnor2 ix7267 (.Y (nx7266), .A0 (nx7264), .A1 (nx3725)) ;
    xnor2 ix7265 (.Y (nx7264), .A0 (nx3977), .A1 (nx7136)) ;
    mux21_ni ix3978 (.Y (nx3977), .A0 (nx3965), .A1 (nx3971), .S0 (nx3967)) ;
    xnor2 ix7137 (.Y (nx7136), .A0 (nx7134), .A1 (nx3983)) ;
    xnor2 ix7135 (.Y (nx7134), .A0 (nx3373), .A1 (nx6992)) ;
    nand02_2x ix3984 (.Y (nx3983), .A0 (input_b[9]), .A1 (input_a[16])) ;
    nand02_2x ix3986 (.Y (nx3985), .A0 (input_b[8]), .A1 (input_a[18])) ;
    xnor2 ix3988 (.Y (nx3987), .A0 (nx3989), .A1 (nx3985)) ;
    xnor2 ix3990 (.Y (nx3989), .A0 (nx3991), .A1 (nx3993)) ;
    mux21_ni ix3992 (.Y (nx3991), .A0 (nx3983), .A1 (nx3977), .S0 (nx7136)) ;
    xnor2 ix3994 (.Y (nx3993), .A0 (nx3995), .A1 (nx3997)) ;
    xnor2 ix3996 (.Y (nx3995), .A0 (nx3369), .A1 (nx3601)) ;
    nand02_2x ix3998 (.Y (nx3997), .A0 (input_b[9]), .A1 (input_a[17])) ;
    xnor2 ix7247 (.Y (nx7246), .A0 (nx7244), .A1 (nx3719)) ;
    xnor2 ix7245 (.Y (nx7244), .A0 (nx4003), .A1 (nx7116)) ;
    mux21_ni ix4004 (.Y (nx4003), .A0 (nx3991), .A1 (nx3997), .S0 (nx3993)) ;
    xnor2 ix7117 (.Y (nx7116), .A0 (nx7114), .A1 (nx4009)) ;
    xnor2 ix7115 (.Y (nx7114), .A0 (nx3367), .A1 (nx6972)) ;
    nand02_2x ix4010 (.Y (nx4009), .A0 (input_b[9]), .A1 (input_a[18])) ;
    nand02_2x ix4012 (.Y (nx4011), .A0 (input_b[8]), .A1 (input_a[20])) ;
    xnor2 ix4014 (.Y (nx4013), .A0 (nx4015), .A1 (nx4011)) ;
    xnor2 ix4016 (.Y (nx4015), .A0 (nx4017), .A1 (nx4019)) ;
    mux21_ni ix4018 (.Y (nx4017), .A0 (nx4009), .A1 (nx4003), .S0 (nx7116)) ;
    xnor2 ix4020 (.Y (nx4019), .A0 (nx4021), .A1 (nx4023)) ;
    xnor2 ix4022 (.Y (nx4021), .A0 (nx3363), .A1 (nx3627)) ;
    nand02_2x ix4024 (.Y (nx4023), .A0 (input_b[9]), .A1 (input_a[19])) ;
    xnor2 ix7227 (.Y (nx7226), .A0 (nx7224), .A1 (nx3713)) ;
    xnor2 ix7225 (.Y (nx7224), .A0 (nx4029), .A1 (nx7096)) ;
    mux21_ni ix4030 (.Y (nx4029), .A0 (nx4017), .A1 (nx4023), .S0 (nx4019)) ;
    xnor2 ix7097 (.Y (nx7096), .A0 (nx7094), .A1 (nx4035)) ;
    xnor2 ix7095 (.Y (nx7094), .A0 (nx3361), .A1 (nx6952)) ;
    nand02_2x ix4036 (.Y (nx4035), .A0 (input_b[9]), .A1 (input_a[20])) ;
    nand02_2x ix4038 (.Y (nx4037), .A0 (input_b[8]), .A1 (input_a[22])) ;
    xnor2 ix4040 (.Y (nx4039), .A0 (nx4041), .A1 (nx4037)) ;
    xnor2 ix4042 (.Y (nx4041), .A0 (nx4043), .A1 (nx4045)) ;
    mux21_ni ix4044 (.Y (nx4043), .A0 (nx4035), .A1 (nx4029), .S0 (nx7096)) ;
    xnor2 ix4046 (.Y (nx4045), .A0 (nx4047), .A1 (nx4049)) ;
    xnor2 ix4048 (.Y (nx4047), .A0 (nx3357), .A1 (nx3653)) ;
    nand02_2x ix4050 (.Y (nx4049), .A0 (input_b[9]), .A1 (input_a[21])) ;
    xnor2 ix4052 (.Y (nx4051), .A0 (input_b[8]), .A1 (nx7204)) ;
    xnor2 ix7205 (.Y (nx7204), .A0 (nx4055), .A1 (nx7076)) ;
    mux21_ni ix4056 (.Y (nx4055), .A0 (nx4043), .A1 (nx4049), .S0 (nx4045)) ;
    xnor2 ix7077 (.Y (nx7076), .A0 (nx7074), .A1 (nx4061)) ;
    xnor2 ix7075 (.Y (nx7074), .A0 (nx3355), .A1 (nx6932)) ;
    nand02_2x ix4062 (.Y (nx4061), .A0 (input_b[9]), .A1 (input_a[22])) ;
    mux21_ni ix4064 (.Y (nx4063), .A0 (nx4065), .A1 (nx5561), .S0 (nx5569)) ;
    mux21_ni ix4066 (.Y (nx4065), .A0 (nx4067), .A1 (nx4423), .S0 (nx7616)) ;
    xnor2 ix4068 (.Y (nx4067), .A0 (nx4069), .A1 (nx4411)) ;
    mux21_ni ix4070 (.Y (nx4069), .A0 (nx4071), .A1 (nx4397), .S0 (nx4399)) ;
    mux21_ni ix4072 (.Y (nx4071), .A0 (nx4073), .A1 (nx4075), .S0 (nx7464)) ;
    nand02_2x ix4074 (.Y (nx4073), .A0 (input_b[6]), .A1 (input_a[21])) ;
    mux21_ni ix4076 (.Y (nx4075), .A0 (nx4077), .A1 (nx4371), .S0 (nx4373)) ;
    mux21_ni ix4078 (.Y (nx4077), .A0 (nx4079), .A1 (nx4081), .S0 (nx7484)) ;
    nand02_2x ix4080 (.Y (nx4079), .A0 (input_b[6]), .A1 (input_a[19])) ;
    mux21_ni ix4082 (.Y (nx4081), .A0 (nx4083), .A1 (nx4345), .S0 (nx4347)) ;
    mux21_ni ix4084 (.Y (nx4083), .A0 (nx4085), .A1 (nx4087), .S0 (nx3888)) ;
    nand02_2x ix4086 (.Y (nx4085), .A0 (input_b[6]), .A1 (input_a[17])) ;
    mux21_ni ix4088 (.Y (nx4087), .A0 (nx4089), .A1 (nx4091), .S0 (nx3290)) ;
    nand02_2x ix4090 (.Y (nx4089), .A0 (input_b[6]), .A1 (input_a[16])) ;
    mux21_ni ix4092 (.Y (nx4091), .A0 (nx4093), .A1 (nx4307), .S0 (nx4309)) ;
    mux21_ni ix4094 (.Y (nx4093), .A0 (nx4095), .A1 (nx4293), .S0 (nx4295)) ;
    mux21_ni ix4096 (.Y (nx4095), .A0 (nx4097), .A1 (nx4279), .S0 (nx4281)) ;
    mux21_ni ix4098 (.Y (nx4097), .A0 (nx4099), .A1 (nx4265), .S0 (nx4267)) ;
    mux21_ni ix4100 (.Y (nx4099), .A0 (nx4101), .A1 (nx4251), .S0 (nx4253)) ;
    mux21_ni ix4102 (.Y (nx4101), .A0 (nx4103), .A1 (nx4237), .S0 (nx4239)) ;
    mux21_ni ix4104 (.Y (nx4103), .A0 (nx4105), .A1 (nx4223), .S0 (nx4225)) ;
    mux21_ni ix4106 (.Y (nx4105), .A0 (nx4107), .A1 (nx4209), .S0 (nx4211)) ;
    mux21_ni ix4108 (.Y (nx4107), .A0 (nx4109), .A1 (nx4195), .S0 (nx4197)) ;
    mux21_ni ix4110 (.Y (nx4109), .A0 (nx4111), .A1 (nx4181), .S0 (nx4183)) ;
    mux21_ni ix4112 (.Y (nx4111), .A0 (nx4113), .A1 (nx4167), .S0 (nx4169)) ;
    mux21_ni ix4114 (.Y (nx4113), .A0 (nx4115), .A1 (nx4151), .S0 (nx4153)) ;
    mux21_ni ix4116 (.Y (nx4115), .A0 (nx4117), .A1 (nx4135), .S0 (nx4137)) ;
    mux21_ni ix4118 (.Y (nx4117), .A0 (nx4119), .A1 (nx4121), .S0 (nx916)) ;
    nand02_2x ix4120 (.Y (nx4119), .A0 (input_b[6]), .A1 (input_a[2])) ;
    xnor2 ix917 (.Y (nx916), .A0 (nx914), .A1 (nx4119)) ;
    inv02 ix4130 (.Y (nx4129), .A (input_b[7])) ;
    inv02 ix4132 (.Y (nx4131), .A (input_b[8])) ;
    aoi22 ix4134 (.Y (nx4133), .A0 (input_b[8]), .A1 (input_a[0]), .B0 (
          input_b[7]), .B1 (input_a[1])) ;
    nand02_2x ix4136 (.Y (nx4135), .A0 (input_b[6]), .A1 (input_a[3])) ;
    xnor2 ix4138 (.Y (nx4137), .A0 (nx4139), .A1 (nx4135)) ;
    xnor2 ix677 (.Y (nx676), .A0 (nx674), .A1 (nx4149)) ;
    aoi22 ix4148 (.Y (nx4147), .A0 (input_b[9]), .A1 (input_a[0]), .B0 (
          input_b[8]), .B1 (input_a[1])) ;
    nand02_2x ix4150 (.Y (nx4149), .A0 (input_b[7]), .A1 (input_a[2])) ;
    nand02_2x ix4152 (.Y (nx4151), .A0 (input_b[6]), .A1 (input_a[4])) ;
    xnor2 ix4154 (.Y (nx4153), .A0 (nx4155), .A1 (nx4151)) ;
    xnor2 ix4156 (.Y (nx4155), .A0 (nx4157), .A1 (nx4161)) ;
    mux21_ni ix4158 (.Y (nx4157), .A0 (nx4149), .A1 (nx4159), .S0 (nx676)) ;
    xnor2 ix4162 (.Y (nx4161), .A0 (nx4163), .A1 (nx4165)) ;
    nand02_2x ix4166 (.Y (nx4165), .A0 (input_b[7]), .A1 (input_a[3])) ;
    nand02_2x ix4168 (.Y (nx4167), .A0 (input_b[6]), .A1 (input_a[5])) ;
    xnor2 ix4170 (.Y (nx4169), .A0 (nx4171), .A1 (nx4167)) ;
    xnor2 ix4172 (.Y (nx4171), .A0 (nx4173), .A1 (nx4175)) ;
    mux21_ni ix4174 (.Y (nx4173), .A0 (nx4157), .A1 (nx4165), .S0 (nx4161)) ;
    xnor2 ix4176 (.Y (nx4175), .A0 (nx4177), .A1 (nx4179)) ;
    xnor2 ix4178 (.Y (nx4177), .A0 (nx3759), .A1 (nx3779)) ;
    nand02_2x ix4180 (.Y (nx4179), .A0 (input_b[7]), .A1 (input_a[4])) ;
    nand02_2x ix4182 (.Y (nx4181), .A0 (input_b[6]), .A1 (input_a[6])) ;
    xnor2 ix4184 (.Y (nx4183), .A0 (nx4185), .A1 (nx4181)) ;
    xnor2 ix4186 (.Y (nx4185), .A0 (nx4187), .A1 (nx4189)) ;
    mux21_ni ix4188 (.Y (nx4187), .A0 (nx4173), .A1 (nx4179), .S0 (nx4175)) ;
    xnor2 ix4190 (.Y (nx4189), .A0 (nx4191), .A1 (nx4193)) ;
    xnor2 ix4192 (.Y (nx4191), .A0 (nx3757), .A1 (nx3795)) ;
    nand02_2x ix4194 (.Y (nx4193), .A0 (input_b[7]), .A1 (input_a[5])) ;
    nand02_2x ix4196 (.Y (nx4195), .A0 (input_b[6]), .A1 (input_a[7])) ;
    xnor2 ix4198 (.Y (nx4197), .A0 (nx4199), .A1 (nx4195)) ;
    xnor2 ix4200 (.Y (nx4199), .A0 (nx4201), .A1 (nx4203)) ;
    mux21_ni ix4202 (.Y (nx4201), .A0 (nx4187), .A1 (nx4193), .S0 (nx4189)) ;
    xnor2 ix4204 (.Y (nx4203), .A0 (nx4205), .A1 (nx4207)) ;
    xnor2 ix4206 (.Y (nx4205), .A0 (nx3755), .A1 (nx3811)) ;
    nand02_2x ix4208 (.Y (nx4207), .A0 (input_b[7]), .A1 (input_a[6])) ;
    nand02_2x ix4210 (.Y (nx4209), .A0 (input_b[6]), .A1 (input_a[8])) ;
    xnor2 ix4212 (.Y (nx4211), .A0 (nx4213), .A1 (nx4209)) ;
    xnor2 ix4214 (.Y (nx4213), .A0 (nx4215), .A1 (nx4217)) ;
    mux21_ni ix4216 (.Y (nx4215), .A0 (nx4201), .A1 (nx4207), .S0 (nx4203)) ;
    xnor2 ix4218 (.Y (nx4217), .A0 (nx4219), .A1 (nx4221)) ;
    xnor2 ix4220 (.Y (nx4219), .A0 (nx3753), .A1 (nx3825)) ;
    nand02_2x ix4222 (.Y (nx4221), .A0 (input_b[7]), .A1 (input_a[7])) ;
    nand02_2x ix4224 (.Y (nx4223), .A0 (input_b[6]), .A1 (input_a[9])) ;
    xnor2 ix4226 (.Y (nx4225), .A0 (nx4227), .A1 (nx4223)) ;
    xnor2 ix4228 (.Y (nx4227), .A0 (nx4229), .A1 (nx4231)) ;
    mux21_ni ix4230 (.Y (nx4229), .A0 (nx4215), .A1 (nx4221), .S0 (nx4217)) ;
    xnor2 ix4232 (.Y (nx4231), .A0 (nx4233), .A1 (nx4235)) ;
    xnor2 ix4234 (.Y (nx4233), .A0 (nx3751), .A1 (nx3839)) ;
    nand02_2x ix4236 (.Y (nx4235), .A0 (input_b[7]), .A1 (input_a[8])) ;
    nand02_2x ix4238 (.Y (nx4237), .A0 (input_b[6]), .A1 (input_a[10])) ;
    xnor2 ix4240 (.Y (nx4239), .A0 (nx4241), .A1 (nx4237)) ;
    xnor2 ix4242 (.Y (nx4241), .A0 (nx4243), .A1 (nx4245)) ;
    mux21_ni ix4244 (.Y (nx4243), .A0 (nx4229), .A1 (nx4235), .S0 (nx4231)) ;
    xnor2 ix4246 (.Y (nx4245), .A0 (nx4247), .A1 (nx4249)) ;
    xnor2 ix4248 (.Y (nx4247), .A0 (nx3749), .A1 (nx3853)) ;
    nand02_2x ix4250 (.Y (nx4249), .A0 (input_b[7]), .A1 (input_a[9])) ;
    nand02_2x ix4252 (.Y (nx4251), .A0 (input_b[6]), .A1 (input_a[11])) ;
    xnor2 ix4254 (.Y (nx4253), .A0 (nx4255), .A1 (nx4251)) ;
    xnor2 ix4256 (.Y (nx4255), .A0 (nx4257), .A1 (nx4259)) ;
    mux21_ni ix4258 (.Y (nx4257), .A0 (nx4243), .A1 (nx4249), .S0 (nx4245)) ;
    xnor2 ix4260 (.Y (nx4259), .A0 (nx4261), .A1 (nx4263)) ;
    xnor2 ix4262 (.Y (nx4261), .A0 (nx3747), .A1 (nx3867)) ;
    nand02_2x ix4264 (.Y (nx4263), .A0 (input_b[7]), .A1 (input_a[10])) ;
    nand02_2x ix4266 (.Y (nx4265), .A0 (input_b[6]), .A1 (input_a[12])) ;
    xnor2 ix4268 (.Y (nx4267), .A0 (nx4269), .A1 (nx4265)) ;
    xnor2 ix4270 (.Y (nx4269), .A0 (nx4271), .A1 (nx4273)) ;
    mux21_ni ix4272 (.Y (nx4271), .A0 (nx4257), .A1 (nx4263), .S0 (nx4259)) ;
    xnor2 ix4274 (.Y (nx4273), .A0 (nx4275), .A1 (nx4277)) ;
    xnor2 ix4276 (.Y (nx4275), .A0 (nx3745), .A1 (nx3881)) ;
    nand02_2x ix4278 (.Y (nx4277), .A0 (input_b[7]), .A1 (input_a[11])) ;
    nand02_2x ix4280 (.Y (nx4279), .A0 (input_b[6]), .A1 (input_a[13])) ;
    xnor2 ix4282 (.Y (nx4281), .A0 (nx4283), .A1 (nx4279)) ;
    xnor2 ix4284 (.Y (nx4283), .A0 (nx4285), .A1 (nx4287)) ;
    mux21_ni ix4286 (.Y (nx4285), .A0 (nx4271), .A1 (nx4277), .S0 (nx4273)) ;
    xnor2 ix4288 (.Y (nx4287), .A0 (nx4289), .A1 (nx4291)) ;
    xnor2 ix4290 (.Y (nx4289), .A0 (nx3743), .A1 (nx3895)) ;
    nand02_2x ix4292 (.Y (nx4291), .A0 (input_b[7]), .A1 (input_a[12])) ;
    nand02_2x ix4294 (.Y (nx4293), .A0 (input_b[6]), .A1 (input_a[14])) ;
    xnor2 ix4296 (.Y (nx4295), .A0 (nx4297), .A1 (nx4293)) ;
    xnor2 ix4298 (.Y (nx4297), .A0 (nx4299), .A1 (nx4301)) ;
    mux21_ni ix4300 (.Y (nx4299), .A0 (nx4285), .A1 (nx4291), .S0 (nx4287)) ;
    xnor2 ix4302 (.Y (nx4301), .A0 (nx4303), .A1 (nx4305)) ;
    xnor2 ix4304 (.Y (nx4303), .A0 (nx3741), .A1 (nx3909)) ;
    nand02_2x ix4306 (.Y (nx4305), .A0 (input_b[7]), .A1 (input_a[13])) ;
    nand02_2x ix4308 (.Y (nx4307), .A0 (input_b[6]), .A1 (input_a[15])) ;
    xnor2 ix4310 (.Y (nx4309), .A0 (nx4311), .A1 (nx4307)) ;
    xnor2 ix4312 (.Y (nx4311), .A0 (nx4313), .A1 (nx4315)) ;
    mux21_ni ix4314 (.Y (nx4313), .A0 (nx4299), .A1 (nx4305), .S0 (nx4301)) ;
    xnor2 ix4316 (.Y (nx4315), .A0 (nx4317), .A1 (nx4319)) ;
    xnor2 ix4318 (.Y (nx4317), .A0 (nx3739), .A1 (nx3923)) ;
    nand02_2x ix4320 (.Y (nx4319), .A0 (input_b[7]), .A1 (input_a[14])) ;
    xnor2 ix3291 (.Y (nx3290), .A0 (nx3286), .A1 (nx4089)) ;
    xnor2 ix3287 (.Y (nx3286), .A0 (nx4325), .A1 (nx3284)) ;
    mux21_ni ix4326 (.Y (nx4325), .A0 (nx4313), .A1 (nx4319), .S0 (nx4315)) ;
    xnor2 ix3285 (.Y (nx3284), .A0 (nx3280), .A1 (nx4331)) ;
    xnor2 ix3281 (.Y (nx3280), .A0 (nx3737), .A1 (nx3278)) ;
    nand02_2x ix4332 (.Y (nx4331), .A0 (input_b[7]), .A1 (input_a[15])) ;
    xnor2 ix3889 (.Y (nx3888), .A0 (nx3884), .A1 (nx4085)) ;
    xnor2 ix3885 (.Y (nx3884), .A0 (nx4337), .A1 (nx3882)) ;
    mux21_ni ix4338 (.Y (nx4337), .A0 (nx4331), .A1 (nx4325), .S0 (nx3284)) ;
    xnor2 ix3883 (.Y (nx3882), .A0 (nx3878), .A1 (nx4343)) ;
    xnor2 ix3879 (.Y (nx3878), .A0 (nx3733), .A1 (nx3876)) ;
    nand02_2x ix4344 (.Y (nx4343), .A0 (input_b[7]), .A1 (input_a[16])) ;
    nand02_2x ix4346 (.Y (nx4345), .A0 (input_b[6]), .A1 (input_a[18])) ;
    xnor2 ix4348 (.Y (nx4347), .A0 (nx4349), .A1 (nx4345)) ;
    xnor2 ix4350 (.Y (nx4349), .A0 (nx4351), .A1 (nx4353)) ;
    mux21_ni ix4352 (.Y (nx4351), .A0 (nx4343), .A1 (nx4337), .S0 (nx3882)) ;
    xnor2 ix4354 (.Y (nx4353), .A0 (nx4355), .A1 (nx4357)) ;
    xnor2 ix4356 (.Y (nx4355), .A0 (nx3729), .A1 (nx3961)) ;
    nand02_2x ix4358 (.Y (nx4357), .A0 (input_b[7]), .A1 (input_a[17])) ;
    xnor2 ix7485 (.Y (nx7484), .A0 (nx7482), .A1 (nx4079)) ;
    xnor2 ix7483 (.Y (nx7482), .A0 (nx4363), .A1 (nx7382)) ;
    mux21_ni ix4364 (.Y (nx4363), .A0 (nx4351), .A1 (nx4357), .S0 (nx4353)) ;
    xnor2 ix7383 (.Y (nx7382), .A0 (nx7380), .A1 (nx4369)) ;
    xnor2 ix7381 (.Y (nx7380), .A0 (nx3727), .A1 (nx7266)) ;
    nand02_2x ix4370 (.Y (nx4369), .A0 (input_b[7]), .A1 (input_a[18])) ;
    nand02_2x ix4372 (.Y (nx4371), .A0 (input_b[6]), .A1 (input_a[20])) ;
    xnor2 ix4374 (.Y (nx4373), .A0 (nx4375), .A1 (nx4371)) ;
    xnor2 ix4376 (.Y (nx4375), .A0 (nx4377), .A1 (nx4379)) ;
    mux21_ni ix4378 (.Y (nx4377), .A0 (nx4369), .A1 (nx4363), .S0 (nx7382)) ;
    xnor2 ix4380 (.Y (nx4379), .A0 (nx4381), .A1 (nx4383)) ;
    xnor2 ix4382 (.Y (nx4381), .A0 (nx3723), .A1 (nx3987)) ;
    nand02_2x ix4384 (.Y (nx4383), .A0 (input_b[7]), .A1 (input_a[19])) ;
    xnor2 ix7465 (.Y (nx7464), .A0 (nx7462), .A1 (nx4073)) ;
    xnor2 ix7463 (.Y (nx7462), .A0 (nx4389), .A1 (nx7362)) ;
    mux21_ni ix4390 (.Y (nx4389), .A0 (nx4377), .A1 (nx4383), .S0 (nx4379)) ;
    xnor2 ix7363 (.Y (nx7362), .A0 (nx7360), .A1 (nx4395)) ;
    xnor2 ix7361 (.Y (nx7360), .A0 (nx3721), .A1 (nx7246)) ;
    nand02_2x ix4396 (.Y (nx4395), .A0 (input_b[7]), .A1 (input_a[20])) ;
    nand02_2x ix4398 (.Y (nx4397), .A0 (input_b[6]), .A1 (input_a[22])) ;
    xnor2 ix4400 (.Y (nx4399), .A0 (nx4401), .A1 (nx4397)) ;
    xnor2 ix4402 (.Y (nx4401), .A0 (nx4403), .A1 (nx4405)) ;
    mux21_ni ix4404 (.Y (nx4403), .A0 (nx4395), .A1 (nx4389), .S0 (nx7362)) ;
    xnor2 ix4406 (.Y (nx4405), .A0 (nx4407), .A1 (nx4409)) ;
    xnor2 ix4408 (.Y (nx4407), .A0 (nx3717), .A1 (nx4013)) ;
    nand02_2x ix4410 (.Y (nx4409), .A0 (input_b[7]), .A1 (input_a[21])) ;
    xnor2 ix4412 (.Y (nx4411), .A0 (input_b[6]), .A1 (nx7442)) ;
    xnor2 ix7443 (.Y (nx7442), .A0 (nx4415), .A1 (nx7342)) ;
    mux21_ni ix4416 (.Y (nx4415), .A0 (nx4403), .A1 (nx4409), .S0 (nx4405)) ;
    xnor2 ix7343 (.Y (nx7342), .A0 (nx7340), .A1 (nx4421)) ;
    xnor2 ix7341 (.Y (nx7340), .A0 (nx3715), .A1 (nx7226)) ;
    nand02_2x ix4422 (.Y (nx4421), .A0 (input_b[7]), .A1 (input_a[22])) ;
    mux21_ni ix7841 (.Y (nx7840), .A0 (nx7692), .A1 (nx7836), .S0 (nx7742)) ;
    mux21_ni ix4430 (.Y (nx4429), .A0 (nx4431), .A1 (nx4757), .S0 (nx4759)) ;
    mux21_ni ix4432 (.Y (nx4431), .A0 (nx4433), .A1 (nx4435), .S0 (nx7646)) ;
    nand02_2x ix4434 (.Y (nx4433), .A0 (input_b[4]), .A1 (input_a[21])) ;
    mux21_ni ix4436 (.Y (nx4435), .A0 (nx4437), .A1 (nx4731), .S0 (nx4733)) ;
    mux21_ni ix4438 (.Y (nx4437), .A0 (nx4439), .A1 (nx4441), .S0 (nx3900)) ;
    nand02_2x ix4440 (.Y (nx4439), .A0 (input_b[4]), .A1 (input_a[19])) ;
    mux21_ni ix4442 (.Y (nx4441), .A0 (nx4443), .A1 (nx4445), .S0 (nx3302)) ;
    nand02_2x ix4444 (.Y (nx4443), .A0 (input_b[4]), .A1 (input_a[18])) ;
    mux21_ni ix4446 (.Y (nx4445), .A0 (nx4447), .A1 (nx4693), .S0 (nx4695)) ;
    mux21_ni ix4448 (.Y (nx4447), .A0 (nx4449), .A1 (nx4679), .S0 (nx4681)) ;
    mux21_ni ix4450 (.Y (nx4449), .A0 (nx4451), .A1 (nx4665), .S0 (nx4667)) ;
    mux21_ni ix4452 (.Y (nx4451), .A0 (nx4453), .A1 (nx4651), .S0 (nx4653)) ;
    mux21_ni ix4454 (.Y (nx4453), .A0 (nx4455), .A1 (nx4637), .S0 (nx4639)) ;
    mux21_ni ix4456 (.Y (nx4455), .A0 (nx4457), .A1 (nx4623), .S0 (nx4625)) ;
    mux21_ni ix4458 (.Y (nx4457), .A0 (nx4459), .A1 (nx4609), .S0 (nx4611)) ;
    mux21_ni ix4460 (.Y (nx4459), .A0 (nx4461), .A1 (nx4595), .S0 (nx4597)) ;
    mux21_ni ix4462 (.Y (nx4461), .A0 (nx4463), .A1 (nx4581), .S0 (nx4583)) ;
    mux21_ni ix4464 (.Y (nx4463), .A0 (nx4465), .A1 (nx4567), .S0 (nx4569)) ;
    mux21_ni ix4466 (.Y (nx4465), .A0 (nx4467), .A1 (nx4553), .S0 (nx4555)) ;
    mux21_ni ix4468 (.Y (nx4467), .A0 (nx4469), .A1 (nx4539), .S0 (nx4541)) ;
    mux21_ni ix4470 (.Y (nx4469), .A0 (nx4471), .A1 (nx4525), .S0 (nx4527)) ;
    mux21_ni ix4472 (.Y (nx4471), .A0 (nx4473), .A1 (nx4509), .S0 (nx4511)) ;
    mux21_ni ix4474 (.Y (nx4473), .A0 (nx4475), .A1 (nx4493), .S0 (nx4495)) ;
    mux21_ni ix4476 (.Y (nx4475), .A0 (nx4477), .A1 (nx4479), .S0 (nx1564)) ;
    nand02_2x ix4478 (.Y (nx4477), .A0 (input_b[4]), .A1 (input_a[2])) ;
    xnor2 ix1565 (.Y (nx1564), .A0 (nx1562), .A1 (nx4477)) ;
    inv02 ix4488 (.Y (nx4487), .A (input_b[5])) ;
    inv02 ix4490 (.Y (nx4489), .A (input_b[6])) ;
    aoi22 ix4492 (.Y (nx4491), .A0 (input_b[6]), .A1 (input_a[0]), .B0 (
          input_b[5]), .B1 (input_a[1])) ;
    nand02_2x ix4494 (.Y (nx4493), .A0 (input_b[4]), .A1 (input_a[3])) ;
    xnor2 ix4496 (.Y (nx4495), .A0 (nx4497), .A1 (nx4493)) ;
    xnor2 ix1213 (.Y (nx1212), .A0 (nx1210), .A1 (nx4507)) ;
    aoi22 ix4506 (.Y (nx4505), .A0 (input_b[7]), .A1 (input_a[0]), .B0 (
          input_b[6]), .B1 (input_a[1])) ;
    nand02_2x ix4508 (.Y (nx4507), .A0 (input_b[5]), .A1 (input_a[2])) ;
    nand02_2x ix4510 (.Y (nx4509), .A0 (input_b[4]), .A1 (input_a[4])) ;
    xnor2 ix4512 (.Y (nx4511), .A0 (nx4513), .A1 (nx4509)) ;
    xnor2 ix4514 (.Y (nx4513), .A0 (nx4515), .A1 (nx4519)) ;
    mux21_ni ix4516 (.Y (nx4515), .A0 (nx4507), .A1 (nx4517), .S0 (nx1212)) ;
    xnor2 ix4520 (.Y (nx4519), .A0 (nx4521), .A1 (nx4523)) ;
    nand02_2x ix4524 (.Y (nx4523), .A0 (input_b[5]), .A1 (input_a[3])) ;
    nand02_2x ix4526 (.Y (nx4525), .A0 (input_b[4]), .A1 (input_a[5])) ;
    xnor2 ix4528 (.Y (nx4527), .A0 (nx4529), .A1 (nx4525)) ;
    xnor2 ix4530 (.Y (nx4529), .A0 (nx4531), .A1 (nx4533)) ;
    mux21_ni ix4532 (.Y (nx4531), .A0 (nx4515), .A1 (nx4523), .S0 (nx4519)) ;
    xnor2 ix4534 (.Y (nx4533), .A0 (nx4535), .A1 (nx4537)) ;
    xnor2 ix4536 (.Y (nx4535), .A0 (nx4117), .A1 (nx4137)) ;
    nand02_2x ix4538 (.Y (nx4537), .A0 (input_b[5]), .A1 (input_a[4])) ;
    nand02_2x ix4540 (.Y (nx4539), .A0 (input_b[4]), .A1 (input_a[6])) ;
    xnor2 ix4542 (.Y (nx4541), .A0 (nx4543), .A1 (nx4539)) ;
    xnor2 ix4544 (.Y (nx4543), .A0 (nx4545), .A1 (nx4547)) ;
    mux21_ni ix4546 (.Y (nx4545), .A0 (nx4531), .A1 (nx4537), .S0 (nx4533)) ;
    xnor2 ix4548 (.Y (nx4547), .A0 (nx4549), .A1 (nx4551)) ;
    xnor2 ix4550 (.Y (nx4549), .A0 (nx4115), .A1 (nx4153)) ;
    nand02_2x ix4552 (.Y (nx4551), .A0 (input_b[5]), .A1 (input_a[5])) ;
    nand02_2x ix4554 (.Y (nx4553), .A0 (input_b[4]), .A1 (input_a[7])) ;
    xnor2 ix4556 (.Y (nx4555), .A0 (nx4557), .A1 (nx4553)) ;
    xnor2 ix4558 (.Y (nx4557), .A0 (nx4559), .A1 (nx4561)) ;
    mux21_ni ix4560 (.Y (nx4559), .A0 (nx4545), .A1 (nx4551), .S0 (nx4547)) ;
    xnor2 ix4562 (.Y (nx4561), .A0 (nx4563), .A1 (nx4565)) ;
    xnor2 ix4564 (.Y (nx4563), .A0 (nx4113), .A1 (nx4169)) ;
    nand02_2x ix4566 (.Y (nx4565), .A0 (input_b[5]), .A1 (input_a[6])) ;
    nand02_2x ix4568 (.Y (nx4567), .A0 (input_b[4]), .A1 (input_a[8])) ;
    xnor2 ix4570 (.Y (nx4569), .A0 (nx4571), .A1 (nx4567)) ;
    xnor2 ix4572 (.Y (nx4571), .A0 (nx4573), .A1 (nx4575)) ;
    mux21_ni ix4574 (.Y (nx4573), .A0 (nx4559), .A1 (nx4565), .S0 (nx4561)) ;
    xnor2 ix4576 (.Y (nx4575), .A0 (nx4577), .A1 (nx4579)) ;
    xnor2 ix4578 (.Y (nx4577), .A0 (nx4111), .A1 (nx4183)) ;
    nand02_2x ix4580 (.Y (nx4579), .A0 (input_b[5]), .A1 (input_a[7])) ;
    nand02_2x ix4582 (.Y (nx4581), .A0 (input_b[4]), .A1 (input_a[9])) ;
    xnor2 ix4584 (.Y (nx4583), .A0 (nx4585), .A1 (nx4581)) ;
    xnor2 ix4586 (.Y (nx4585), .A0 (nx4587), .A1 (nx4589)) ;
    mux21_ni ix4588 (.Y (nx4587), .A0 (nx4573), .A1 (nx4579), .S0 (nx4575)) ;
    xnor2 ix4590 (.Y (nx4589), .A0 (nx4591), .A1 (nx4593)) ;
    xnor2 ix4592 (.Y (nx4591), .A0 (nx4109), .A1 (nx4197)) ;
    nand02_2x ix4594 (.Y (nx4593), .A0 (input_b[5]), .A1 (input_a[8])) ;
    nand02_2x ix4596 (.Y (nx4595), .A0 (input_b[4]), .A1 (input_a[10])) ;
    xnor2 ix4598 (.Y (nx4597), .A0 (nx4599), .A1 (nx4595)) ;
    xnor2 ix4600 (.Y (nx4599), .A0 (nx4601), .A1 (nx4603)) ;
    mux21_ni ix4602 (.Y (nx4601), .A0 (nx4587), .A1 (nx4593), .S0 (nx4589)) ;
    xnor2 ix4604 (.Y (nx4603), .A0 (nx4605), .A1 (nx4607)) ;
    xnor2 ix4606 (.Y (nx4605), .A0 (nx4107), .A1 (nx4211)) ;
    nand02_2x ix4608 (.Y (nx4607), .A0 (input_b[5]), .A1 (input_a[9])) ;
    nand02_2x ix4610 (.Y (nx4609), .A0 (input_b[4]), .A1 (input_a[11])) ;
    xnor2 ix4612 (.Y (nx4611), .A0 (nx4613), .A1 (nx4609)) ;
    xnor2 ix4614 (.Y (nx4613), .A0 (nx4615), .A1 (nx4617)) ;
    mux21_ni ix4616 (.Y (nx4615), .A0 (nx4601), .A1 (nx4607), .S0 (nx4603)) ;
    xnor2 ix4618 (.Y (nx4617), .A0 (nx4619), .A1 (nx4621)) ;
    xnor2 ix4620 (.Y (nx4619), .A0 (nx4105), .A1 (nx4225)) ;
    nand02_2x ix4622 (.Y (nx4621), .A0 (input_b[5]), .A1 (input_a[10])) ;
    nand02_2x ix4624 (.Y (nx4623), .A0 (input_b[4]), .A1 (input_a[12])) ;
    xnor2 ix4626 (.Y (nx4625), .A0 (nx4627), .A1 (nx4623)) ;
    xnor2 ix4628 (.Y (nx4627), .A0 (nx4629), .A1 (nx4631)) ;
    mux21_ni ix4630 (.Y (nx4629), .A0 (nx4615), .A1 (nx4621), .S0 (nx4617)) ;
    xnor2 ix4632 (.Y (nx4631), .A0 (nx4633), .A1 (nx4635)) ;
    xnor2 ix4634 (.Y (nx4633), .A0 (nx4103), .A1 (nx4239)) ;
    nand02_2x ix4636 (.Y (nx4635), .A0 (input_b[5]), .A1 (input_a[11])) ;
    nand02_2x ix4638 (.Y (nx4637), .A0 (input_b[4]), .A1 (input_a[13])) ;
    xnor2 ix4640 (.Y (nx4639), .A0 (nx4641), .A1 (nx4637)) ;
    xnor2 ix4642 (.Y (nx4641), .A0 (nx4643), .A1 (nx4645)) ;
    mux21_ni ix4644 (.Y (nx4643), .A0 (nx4629), .A1 (nx4635), .S0 (nx4631)) ;
    xnor2 ix4646 (.Y (nx4645), .A0 (nx4647), .A1 (nx4649)) ;
    xnor2 ix4648 (.Y (nx4647), .A0 (nx4101), .A1 (nx4253)) ;
    nand02_2x ix4650 (.Y (nx4649), .A0 (input_b[5]), .A1 (input_a[12])) ;
    nand02_2x ix4652 (.Y (nx4651), .A0 (input_b[4]), .A1 (input_a[14])) ;
    xnor2 ix4654 (.Y (nx4653), .A0 (nx4655), .A1 (nx4651)) ;
    xnor2 ix4656 (.Y (nx4655), .A0 (nx4657), .A1 (nx4659)) ;
    mux21_ni ix4658 (.Y (nx4657), .A0 (nx4643), .A1 (nx4649), .S0 (nx4645)) ;
    xnor2 ix4660 (.Y (nx4659), .A0 (nx4661), .A1 (nx4663)) ;
    xnor2 ix4662 (.Y (nx4661), .A0 (nx4099), .A1 (nx4267)) ;
    nand02_2x ix4664 (.Y (nx4663), .A0 (input_b[5]), .A1 (input_a[13])) ;
    nand02_2x ix4666 (.Y (nx4665), .A0 (input_b[4]), .A1 (input_a[15])) ;
    xnor2 ix4668 (.Y (nx4667), .A0 (nx4669), .A1 (nx4665)) ;
    xnor2 ix4670 (.Y (nx4669), .A0 (nx4671), .A1 (nx4673)) ;
    mux21_ni ix4672 (.Y (nx4671), .A0 (nx4657), .A1 (nx4663), .S0 (nx4659)) ;
    xnor2 ix4674 (.Y (nx4673), .A0 (nx4675), .A1 (nx4677)) ;
    xnor2 ix4676 (.Y (nx4675), .A0 (nx4097), .A1 (nx4281)) ;
    nand02_2x ix4678 (.Y (nx4677), .A0 (input_b[5]), .A1 (input_a[14])) ;
    nand02_2x ix4680 (.Y (nx4679), .A0 (input_b[4]), .A1 (input_a[16])) ;
    xnor2 ix4682 (.Y (nx4681), .A0 (nx4683), .A1 (nx4679)) ;
    xnor2 ix4684 (.Y (nx4683), .A0 (nx4685), .A1 (nx4687)) ;
    mux21_ni ix4686 (.Y (nx4685), .A0 (nx4671), .A1 (nx4677), .S0 (nx4673)) ;
    xnor2 ix4688 (.Y (nx4687), .A0 (nx4689), .A1 (nx4691)) ;
    xnor2 ix4690 (.Y (nx4689), .A0 (nx4095), .A1 (nx4295)) ;
    nand02_2x ix4692 (.Y (nx4691), .A0 (input_b[5]), .A1 (input_a[15])) ;
    nand02_2x ix4694 (.Y (nx4693), .A0 (input_b[4]), .A1 (input_a[17])) ;
    xnor2 ix4696 (.Y (nx4695), .A0 (nx4697), .A1 (nx4693)) ;
    xnor2 ix4698 (.Y (nx4697), .A0 (nx4699), .A1 (nx4701)) ;
    mux21_ni ix4700 (.Y (nx4699), .A0 (nx4685), .A1 (nx4691), .S0 (nx4687)) ;
    xnor2 ix4702 (.Y (nx4701), .A0 (nx4703), .A1 (nx4705)) ;
    xnor2 ix4704 (.Y (nx4703), .A0 (nx4093), .A1 (nx4309)) ;
    nand02_2x ix4706 (.Y (nx4705), .A0 (input_b[5]), .A1 (input_a[16])) ;
    xnor2 ix3303 (.Y (nx3302), .A0 (nx3298), .A1 (nx4443)) ;
    xnor2 ix3299 (.Y (nx3298), .A0 (nx4711), .A1 (nx3296)) ;
    mux21_ni ix4712 (.Y (nx4711), .A0 (nx4699), .A1 (nx4705), .S0 (nx4701)) ;
    xnor2 ix3297 (.Y (nx3296), .A0 (nx3292), .A1 (nx4717)) ;
    xnor2 ix3293 (.Y (nx3292), .A0 (nx4091), .A1 (nx3290)) ;
    nand02_2x ix4718 (.Y (nx4717), .A0 (input_b[5]), .A1 (input_a[17])) ;
    xnor2 ix3901 (.Y (nx3900), .A0 (nx3896), .A1 (nx4439)) ;
    xnor2 ix3897 (.Y (nx3896), .A0 (nx4723), .A1 (nx3894)) ;
    mux21_ni ix4724 (.Y (nx4723), .A0 (nx4717), .A1 (nx4711), .S0 (nx3296)) ;
    xnor2 ix3895 (.Y (nx3894), .A0 (nx3890), .A1 (nx4729)) ;
    xnor2 ix3891 (.Y (nx3890), .A0 (nx4087), .A1 (nx3888)) ;
    nand02_2x ix4730 (.Y (nx4729), .A0 (input_b[5]), .A1 (input_a[18])) ;
    nand02_2x ix4732 (.Y (nx4731), .A0 (input_b[4]), .A1 (input_a[20])) ;
    xnor2 ix4734 (.Y (nx4733), .A0 (nx4735), .A1 (nx4731)) ;
    xnor2 ix4736 (.Y (nx4735), .A0 (nx4737), .A1 (nx4739)) ;
    mux21_ni ix4738 (.Y (nx4737), .A0 (nx4729), .A1 (nx4723), .S0 (nx3894)) ;
    xnor2 ix4740 (.Y (nx4739), .A0 (nx4741), .A1 (nx4743)) ;
    xnor2 ix4742 (.Y (nx4741), .A0 (nx4083), .A1 (nx4347)) ;
    nand02_2x ix4744 (.Y (nx4743), .A0 (input_b[5]), .A1 (input_a[19])) ;
    xnor2 ix7647 (.Y (nx7646), .A0 (nx7644), .A1 (nx4433)) ;
    xnor2 ix7645 (.Y (nx7644), .A0 (nx4749), .A1 (nx7572)) ;
    mux21_ni ix4750 (.Y (nx4749), .A0 (nx4737), .A1 (nx4743), .S0 (nx4739)) ;
    xnor2 ix7573 (.Y (nx7572), .A0 (nx7570), .A1 (nx4755)) ;
    xnor2 ix7571 (.Y (nx7570), .A0 (nx4081), .A1 (nx7484)) ;
    nand02_2x ix4756 (.Y (nx4755), .A0 (input_b[5]), .A1 (input_a[20])) ;
    nand02_2x ix4758 (.Y (nx4757), .A0 (input_b[4]), .A1 (input_a[22])) ;
    xnor2 ix4760 (.Y (nx4759), .A0 (nx4761), .A1 (nx4757)) ;
    xnor2 ix4762 (.Y (nx4761), .A0 (nx4763), .A1 (nx4765)) ;
    mux21_ni ix4764 (.Y (nx4763), .A0 (nx4755), .A1 (nx4749), .S0 (nx7572)) ;
    xnor2 ix4766 (.Y (nx4765), .A0 (nx4767), .A1 (nx4769)) ;
    xnor2 ix4768 (.Y (nx4767), .A0 (nx4077), .A1 (nx4373)) ;
    nand02_2x ix4770 (.Y (nx4769), .A0 (input_b[5]), .A1 (input_a[21])) ;
    xnor2 ix4772 (.Y (nx4771), .A0 (input_b[4]), .A1 (nx7624)) ;
    xnor2 ix7625 (.Y (nx7624), .A0 (nx4775), .A1 (nx7552)) ;
    mux21_ni ix4776 (.Y (nx4775), .A0 (nx4763), .A1 (nx4769), .S0 (nx4765)) ;
    xnor2 ix7553 (.Y (nx7552), .A0 (nx7550), .A1 (nx4781)) ;
    xnor2 ix7551 (.Y (nx7550), .A0 (nx4075), .A1 (nx7464)) ;
    nand02_2x ix4782 (.Y (nx4781), .A0 (input_b[5]), .A1 (input_a[22])) ;
    mux21_ni ix7837 (.Y (nx7836), .A0 (nx7832), .A1 (nx7748), .S0 (nx5527)) ;
    xnor2 ix4788 (.Y (nx4787), .A0 (nx4789), .A1 (nx5131)) ;
    mux21_ni ix4790 (.Y (nx4789), .A0 (nx4791), .A1 (nx5117), .S0 (nx5119)) ;
    mux21_ni ix4792 (.Y (nx4791), .A0 (nx4793), .A1 (nx4795), .S0 (nx3912)) ;
    nand02_2x ix4794 (.Y (nx4793), .A0 (input_b[2]), .A1 (input_a[21])) ;
    mux21_ni ix4796 (.Y (nx4795), .A0 (nx4797), .A1 (nx4799), .S0 (nx3314)) ;
    nand02_2x ix4798 (.Y (nx4797), .A0 (input_b[2]), .A1 (input_a[20])) ;
    mux21_ni ix4800 (.Y (nx4799), .A0 (nx4801), .A1 (nx5079), .S0 (nx5081)) ;
    mux21_ni ix4802 (.Y (nx4801), .A0 (nx4803), .A1 (nx5065), .S0 (nx5067)) ;
    mux21_ni ix4804 (.Y (nx4803), .A0 (nx4805), .A1 (nx5051), .S0 (nx5053)) ;
    mux21_ni ix4806 (.Y (nx4805), .A0 (nx4807), .A1 (nx5037), .S0 (nx5039)) ;
    mux21_ni ix4808 (.Y (nx4807), .A0 (nx4809), .A1 (nx5023), .S0 (nx5025)) ;
    mux21_ni ix4810 (.Y (nx4809), .A0 (nx4811), .A1 (nx5009), .S0 (nx5011)) ;
    mux21_ni ix4812 (.Y (nx4811), .A0 (nx4813), .A1 (nx4995), .S0 (nx4997)) ;
    mux21_ni ix4814 (.Y (nx4813), .A0 (nx4815), .A1 (nx4981), .S0 (nx4983)) ;
    mux21_ni ix4816 (.Y (nx4815), .A0 (nx4817), .A1 (nx4967), .S0 (nx4969)) ;
    mux21_ni ix4818 (.Y (nx4817), .A0 (nx4819), .A1 (nx4953), .S0 (nx4955)) ;
    mux21_ni ix4820 (.Y (nx4819), .A0 (nx4821), .A1 (nx4939), .S0 (nx4941)) ;
    mux21_ni ix4822 (.Y (nx4821), .A0 (nx4823), .A1 (nx4925), .S0 (nx4927)) ;
    mux21_ni ix4824 (.Y (nx4823), .A0 (nx4825), .A1 (nx4911), .S0 (nx4913)) ;
    mux21_ni ix4826 (.Y (nx4825), .A0 (nx4827), .A1 (nx4897), .S0 (nx4899)) ;
    mux21_ni ix4828 (.Y (nx4827), .A0 (nx4829), .A1 (nx4883), .S0 (nx4885)) ;
    mux21_ni ix4830 (.Y (nx4829), .A0 (nx4831), .A1 (nx4867), .S0 (nx4869)) ;
    mux21_ni ix4832 (.Y (nx4831), .A0 (nx4833), .A1 (nx4851), .S0 (nx4853)) ;
    mux21_ni ix4834 (.Y (nx4833), .A0 (nx4835), .A1 (nx4837), .S0 (nx2436)) ;
    nand02_2x ix4836 (.Y (nx4835), .A0 (input_b[2]), .A1 (input_a[2])) ;
    xnor2 ix2437 (.Y (nx2436), .A0 (nx2434), .A1 (nx4835)) ;
    inv02 ix4846 (.Y (nx4845), .A (input_b[3])) ;
    inv02 ix4848 (.Y (nx4847), .A (input_b[4])) ;
    aoi22 ix4850 (.Y (nx4849), .A0 (input_b[4]), .A1 (input_a[0]), .B0 (
          input_b[3]), .B1 (input_a[1])) ;
    nand02_2x ix4852 (.Y (nx4851), .A0 (input_b[2]), .A1 (input_a[3])) ;
    xnor2 ix4854 (.Y (nx4853), .A0 (nx4855), .A1 (nx4851)) ;
    xnor2 ix1973 (.Y (nx1972), .A0 (nx1970), .A1 (nx4865)) ;
    aoi22 ix4864 (.Y (nx4863), .A0 (input_b[5]), .A1 (input_a[0]), .B0 (
          input_b[4]), .B1 (input_a[1])) ;
    nand02_2x ix4866 (.Y (nx4865), .A0 (input_b[3]), .A1 (input_a[2])) ;
    nand02_2x ix4868 (.Y (nx4867), .A0 (input_b[2]), .A1 (input_a[4])) ;
    xnor2 ix4870 (.Y (nx4869), .A0 (nx4871), .A1 (nx4867)) ;
    xnor2 ix4872 (.Y (nx4871), .A0 (nx4873), .A1 (nx4877)) ;
    mux21_ni ix4874 (.Y (nx4873), .A0 (nx4865), .A1 (nx4875), .S0 (nx1972)) ;
    xnor2 ix4878 (.Y (nx4877), .A0 (nx4879), .A1 (nx4881)) ;
    nand02_2x ix4882 (.Y (nx4881), .A0 (input_b[3]), .A1 (input_a[3])) ;
    nand02_2x ix4884 (.Y (nx4883), .A0 (input_b[2]), .A1 (input_a[5])) ;
    xnor2 ix4886 (.Y (nx4885), .A0 (nx4887), .A1 (nx4883)) ;
    xnor2 ix4888 (.Y (nx4887), .A0 (nx4889), .A1 (nx4891)) ;
    mux21_ni ix4890 (.Y (nx4889), .A0 (nx4873), .A1 (nx4881), .S0 (nx4877)) ;
    xnor2 ix4892 (.Y (nx4891), .A0 (nx4893), .A1 (nx4895)) ;
    xnor2 ix4894 (.Y (nx4893), .A0 (nx4475), .A1 (nx4495)) ;
    nand02_2x ix4896 (.Y (nx4895), .A0 (input_b[3]), .A1 (input_a[4])) ;
    nand02_2x ix4898 (.Y (nx4897), .A0 (input_b[2]), .A1 (input_a[6])) ;
    xnor2 ix4900 (.Y (nx4899), .A0 (nx4901), .A1 (nx4897)) ;
    xnor2 ix4902 (.Y (nx4901), .A0 (nx4903), .A1 (nx4905)) ;
    mux21_ni ix4904 (.Y (nx4903), .A0 (nx4889), .A1 (nx4895), .S0 (nx4891)) ;
    xnor2 ix4906 (.Y (nx4905), .A0 (nx4907), .A1 (nx4909)) ;
    xnor2 ix4908 (.Y (nx4907), .A0 (nx4473), .A1 (nx4511)) ;
    nand02_2x ix4910 (.Y (nx4909), .A0 (input_b[3]), .A1 (input_a[5])) ;
    nand02_2x ix4912 (.Y (nx4911), .A0 (input_b[2]), .A1 (input_a[7])) ;
    xnor2 ix4914 (.Y (nx4913), .A0 (nx4915), .A1 (nx4911)) ;
    xnor2 ix4916 (.Y (nx4915), .A0 (nx4917), .A1 (nx4919)) ;
    mux21_ni ix4918 (.Y (nx4917), .A0 (nx4903), .A1 (nx4909), .S0 (nx4905)) ;
    xnor2 ix4920 (.Y (nx4919), .A0 (nx4921), .A1 (nx4923)) ;
    xnor2 ix4922 (.Y (nx4921), .A0 (nx4471), .A1 (nx4527)) ;
    nand02_2x ix4924 (.Y (nx4923), .A0 (input_b[3]), .A1 (input_a[6])) ;
    nand02_2x ix4926 (.Y (nx4925), .A0 (input_b[2]), .A1 (input_a[8])) ;
    xnor2 ix4928 (.Y (nx4927), .A0 (nx4929), .A1 (nx4925)) ;
    xnor2 ix4930 (.Y (nx4929), .A0 (nx4931), .A1 (nx4933)) ;
    mux21_ni ix4932 (.Y (nx4931), .A0 (nx4917), .A1 (nx4923), .S0 (nx4919)) ;
    xnor2 ix4934 (.Y (nx4933), .A0 (nx4935), .A1 (nx4937)) ;
    xnor2 ix4936 (.Y (nx4935), .A0 (nx4469), .A1 (nx4541)) ;
    nand02_2x ix4938 (.Y (nx4937), .A0 (input_b[3]), .A1 (input_a[7])) ;
    nand02_2x ix4940 (.Y (nx4939), .A0 (input_b[2]), .A1 (input_a[9])) ;
    xnor2 ix4942 (.Y (nx4941), .A0 (nx4943), .A1 (nx4939)) ;
    xnor2 ix4944 (.Y (nx4943), .A0 (nx4945), .A1 (nx4947)) ;
    mux21_ni ix4946 (.Y (nx4945), .A0 (nx4931), .A1 (nx4937), .S0 (nx4933)) ;
    xnor2 ix4948 (.Y (nx4947), .A0 (nx4949), .A1 (nx4951)) ;
    xnor2 ix4950 (.Y (nx4949), .A0 (nx4467), .A1 (nx4555)) ;
    nand02_2x ix4952 (.Y (nx4951), .A0 (input_b[3]), .A1 (input_a[8])) ;
    nand02_2x ix4954 (.Y (nx4953), .A0 (input_b[2]), .A1 (input_a[10])) ;
    xnor2 ix4956 (.Y (nx4955), .A0 (nx4957), .A1 (nx4953)) ;
    xnor2 ix4958 (.Y (nx4957), .A0 (nx4959), .A1 (nx4961)) ;
    mux21_ni ix4960 (.Y (nx4959), .A0 (nx4945), .A1 (nx4951), .S0 (nx4947)) ;
    xnor2 ix4962 (.Y (nx4961), .A0 (nx4963), .A1 (nx4965)) ;
    xnor2 ix4964 (.Y (nx4963), .A0 (nx4465), .A1 (nx4569)) ;
    nand02_2x ix4966 (.Y (nx4965), .A0 (input_b[3]), .A1 (input_a[9])) ;
    nand02_2x ix4968 (.Y (nx4967), .A0 (input_b[2]), .A1 (input_a[11])) ;
    xnor2 ix4970 (.Y (nx4969), .A0 (nx4971), .A1 (nx4967)) ;
    xnor2 ix4972 (.Y (nx4971), .A0 (nx4973), .A1 (nx4975)) ;
    mux21_ni ix4974 (.Y (nx4973), .A0 (nx4959), .A1 (nx4965), .S0 (nx4961)) ;
    xnor2 ix4976 (.Y (nx4975), .A0 (nx4977), .A1 (nx4979)) ;
    xnor2 ix4978 (.Y (nx4977), .A0 (nx4463), .A1 (nx4583)) ;
    nand02_2x ix4980 (.Y (nx4979), .A0 (input_b[3]), .A1 (input_a[10])) ;
    nand02_2x ix4982 (.Y (nx4981), .A0 (input_b[2]), .A1 (input_a[12])) ;
    xnor2 ix4984 (.Y (nx4983), .A0 (nx4985), .A1 (nx4981)) ;
    xnor2 ix4986 (.Y (nx4985), .A0 (nx4987), .A1 (nx4989)) ;
    mux21_ni ix4988 (.Y (nx4987), .A0 (nx4973), .A1 (nx4979), .S0 (nx4975)) ;
    xnor2 ix4990 (.Y (nx4989), .A0 (nx4991), .A1 (nx4993)) ;
    xnor2 ix4992 (.Y (nx4991), .A0 (nx4461), .A1 (nx4597)) ;
    nand02_2x ix4994 (.Y (nx4993), .A0 (input_b[3]), .A1 (input_a[11])) ;
    nand02_2x ix4996 (.Y (nx4995), .A0 (input_b[2]), .A1 (input_a[13])) ;
    xnor2 ix4998 (.Y (nx4997), .A0 (nx4999), .A1 (nx4995)) ;
    xnor2 ix5000 (.Y (nx4999), .A0 (nx5001), .A1 (nx5003)) ;
    mux21_ni ix5002 (.Y (nx5001), .A0 (nx4987), .A1 (nx4993), .S0 (nx4989)) ;
    xnor2 ix5004 (.Y (nx5003), .A0 (nx5005), .A1 (nx5007)) ;
    xnor2 ix5006 (.Y (nx5005), .A0 (nx4459), .A1 (nx4611)) ;
    nand02_2x ix5008 (.Y (nx5007), .A0 (input_b[3]), .A1 (input_a[12])) ;
    nand02_2x ix5010 (.Y (nx5009), .A0 (input_b[2]), .A1 (input_a[14])) ;
    xnor2 ix5012 (.Y (nx5011), .A0 (nx5013), .A1 (nx5009)) ;
    xnor2 ix5014 (.Y (nx5013), .A0 (nx5015), .A1 (nx5017)) ;
    mux21_ni ix5016 (.Y (nx5015), .A0 (nx5001), .A1 (nx5007), .S0 (nx5003)) ;
    xnor2 ix5018 (.Y (nx5017), .A0 (nx5019), .A1 (nx5021)) ;
    xnor2 ix5020 (.Y (nx5019), .A0 (nx4457), .A1 (nx4625)) ;
    nand02_2x ix5022 (.Y (nx5021), .A0 (input_b[3]), .A1 (input_a[13])) ;
    nand02_2x ix5024 (.Y (nx5023), .A0 (input_b[2]), .A1 (input_a[15])) ;
    xnor2 ix5026 (.Y (nx5025), .A0 (nx5027), .A1 (nx5023)) ;
    xnor2 ix5028 (.Y (nx5027), .A0 (nx5029), .A1 (nx5031)) ;
    mux21_ni ix5030 (.Y (nx5029), .A0 (nx5015), .A1 (nx5021), .S0 (nx5017)) ;
    xnor2 ix5032 (.Y (nx5031), .A0 (nx5033), .A1 (nx5035)) ;
    xnor2 ix5034 (.Y (nx5033), .A0 (nx4455), .A1 (nx4639)) ;
    nand02_2x ix5036 (.Y (nx5035), .A0 (input_b[3]), .A1 (input_a[14])) ;
    nand02_2x ix5038 (.Y (nx5037), .A0 (input_b[2]), .A1 (input_a[16])) ;
    xnor2 ix5040 (.Y (nx5039), .A0 (nx5041), .A1 (nx5037)) ;
    xnor2 ix5042 (.Y (nx5041), .A0 (nx5043), .A1 (nx5045)) ;
    mux21_ni ix5044 (.Y (nx5043), .A0 (nx5029), .A1 (nx5035), .S0 (nx5031)) ;
    xnor2 ix5046 (.Y (nx5045), .A0 (nx5047), .A1 (nx5049)) ;
    xnor2 ix5048 (.Y (nx5047), .A0 (nx4453), .A1 (nx4653)) ;
    nand02_2x ix5050 (.Y (nx5049), .A0 (input_b[3]), .A1 (input_a[15])) ;
    nand02_2x ix5052 (.Y (nx5051), .A0 (input_b[2]), .A1 (input_a[17])) ;
    xnor2 ix5054 (.Y (nx5053), .A0 (nx5055), .A1 (nx5051)) ;
    xnor2 ix5056 (.Y (nx5055), .A0 (nx5057), .A1 (nx5059)) ;
    mux21_ni ix5058 (.Y (nx5057), .A0 (nx5043), .A1 (nx5049), .S0 (nx5045)) ;
    xnor2 ix5060 (.Y (nx5059), .A0 (nx5061), .A1 (nx5063)) ;
    xnor2 ix5062 (.Y (nx5061), .A0 (nx4451), .A1 (nx4667)) ;
    nand02_2x ix5064 (.Y (nx5063), .A0 (input_b[3]), .A1 (input_a[16])) ;
    nand02_2x ix5066 (.Y (nx5065), .A0 (input_b[2]), .A1 (input_a[18])) ;
    xnor2 ix5068 (.Y (nx5067), .A0 (nx5069), .A1 (nx5065)) ;
    xnor2 ix5070 (.Y (nx5069), .A0 (nx5071), .A1 (nx5073)) ;
    mux21_ni ix5072 (.Y (nx5071), .A0 (nx5057), .A1 (nx5063), .S0 (nx5059)) ;
    xnor2 ix5074 (.Y (nx5073), .A0 (nx5075), .A1 (nx5077)) ;
    xnor2 ix5076 (.Y (nx5075), .A0 (nx4449), .A1 (nx4681)) ;
    nand02_2x ix5078 (.Y (nx5077), .A0 (input_b[3]), .A1 (input_a[17])) ;
    nand02_2x ix5080 (.Y (nx5079), .A0 (input_b[2]), .A1 (input_a[19])) ;
    xnor2 ix5082 (.Y (nx5081), .A0 (nx5083), .A1 (nx5079)) ;
    xnor2 ix5084 (.Y (nx5083), .A0 (nx5085), .A1 (nx5087)) ;
    mux21_ni ix5086 (.Y (nx5085), .A0 (nx5071), .A1 (nx5077), .S0 (nx5073)) ;
    xnor2 ix5088 (.Y (nx5087), .A0 (nx5089), .A1 (nx5091)) ;
    xnor2 ix5090 (.Y (nx5089), .A0 (nx4447), .A1 (nx4695)) ;
    nand02_2x ix5092 (.Y (nx5091), .A0 (input_b[3]), .A1 (input_a[18])) ;
    xnor2 ix3315 (.Y (nx3314), .A0 (nx3310), .A1 (nx4797)) ;
    xnor2 ix3311 (.Y (nx3310), .A0 (nx5097), .A1 (nx3308)) ;
    mux21_ni ix5098 (.Y (nx5097), .A0 (nx5085), .A1 (nx5091), .S0 (nx5087)) ;
    xnor2 ix3309 (.Y (nx3308), .A0 (nx3304), .A1 (nx5103)) ;
    xnor2 ix3305 (.Y (nx3304), .A0 (nx4445), .A1 (nx3302)) ;
    nand02_2x ix5104 (.Y (nx5103), .A0 (input_b[3]), .A1 (input_a[19])) ;
    xnor2 ix3913 (.Y (nx3912), .A0 (nx3908), .A1 (nx4793)) ;
    xnor2 ix3909 (.Y (nx3908), .A0 (nx5109), .A1 (nx3906)) ;
    mux21_ni ix5110 (.Y (nx5109), .A0 (nx5103), .A1 (nx5097), .S0 (nx3308)) ;
    xnor2 ix3907 (.Y (nx3906), .A0 (nx3902), .A1 (nx5115)) ;
    xnor2 ix3903 (.Y (nx3902), .A0 (nx4441), .A1 (nx3900)) ;
    nand02_2x ix5116 (.Y (nx5115), .A0 (input_b[3]), .A1 (input_a[20])) ;
    nand02_2x ix5118 (.Y (nx5117), .A0 (input_b[2]), .A1 (input_a[22])) ;
    xnor2 ix5120 (.Y (nx5119), .A0 (nx5121), .A1 (nx5117)) ;
    xnor2 ix5122 (.Y (nx5121), .A0 (nx5123), .A1 (nx5125)) ;
    mux21_ni ix5124 (.Y (nx5123), .A0 (nx5115), .A1 (nx5109), .S0 (nx3906)) ;
    xnor2 ix5126 (.Y (nx5125), .A0 (nx5127), .A1 (nx5129)) ;
    xnor2 ix5128 (.Y (nx5127), .A0 (nx4437), .A1 (nx4733)) ;
    nand02_2x ix5130 (.Y (nx5129), .A0 (input_b[3]), .A1 (input_a[21])) ;
    xnor2 ix5132 (.Y (nx5131), .A0 (input_b[2]), .A1 (nx7750)) ;
    xnor2 ix7751 (.Y (nx7750), .A0 (nx5135), .A1 (nx7706)) ;
    mux21_ni ix5136 (.Y (nx5135), .A0 (nx5123), .A1 (nx5129), .S0 (nx5125)) ;
    xnor2 ix7707 (.Y (nx7706), .A0 (nx7704), .A1 (nx5141)) ;
    xnor2 ix7705 (.Y (nx7704), .A0 (nx4435), .A1 (nx7646)) ;
    nand02_2x ix5142 (.Y (nx5141), .A0 (input_b[3]), .A1 (input_a[22])) ;
    nand02_2x ix5144 (.Y (nx5143), .A0 (nx7824), .A1 (nx7826)) ;
    oai22 ix7825 (.Y (nx7824), .A0 (nx5147), .A1 (nx5323), .B0 (nx5325), .B1 (
          nx5501)) ;
    mux21_ni ix5150 (.Y (nx5149), .A0 (nx5151), .A1 (nx5153), .S0 (nx3320)) ;
    nand02_2x ix5152 (.Y (nx5151), .A0 (input_b[1]), .A1 (input_a[21])) ;
    mux21_ni ix5154 (.Y (nx5153), .A0 (nx5155), .A1 (nx5307), .S0 (nx5309)) ;
    mux21_ni ix5156 (.Y (nx5155), .A0 (nx5157), .A1 (nx5301), .S0 (nx5303)) ;
    mux21_ni ix5158 (.Y (nx5157), .A0 (nx5159), .A1 (nx5295), .S0 (nx5297)) ;
    mux21_ni ix5160 (.Y (nx5159), .A0 (nx5161), .A1 (nx5289), .S0 (nx5291)) ;
    mux21_ni ix5162 (.Y (nx5161), .A0 (nx5163), .A1 (nx5283), .S0 (nx5285)) ;
    mux21_ni ix5164 (.Y (nx5163), .A0 (nx5165), .A1 (nx5277), .S0 (nx5279)) ;
    mux21_ni ix5166 (.Y (nx5165), .A0 (nx5167), .A1 (nx5271), .S0 (nx5273)) ;
    mux21_ni ix5168 (.Y (nx5167), .A0 (nx5169), .A1 (nx5265), .S0 (nx5267)) ;
    mux21_ni ix5170 (.Y (nx5169), .A0 (nx5171), .A1 (nx5259), .S0 (nx5261)) ;
    mux21_ni ix5172 (.Y (nx5171), .A0 (nx5173), .A1 (nx5253), .S0 (nx5255)) ;
    mux21_ni ix5174 (.Y (nx5173), .A0 (nx5175), .A1 (nx5247), .S0 (nx5249)) ;
    mux21_ni ix5176 (.Y (nx5175), .A0 (nx5177), .A1 (nx5241), .S0 (nx5243)) ;
    mux21_ni ix5178 (.Y (nx5177), .A0 (nx5179), .A1 (nx5235), .S0 (nx5237)) ;
    mux21_ni ix5180 (.Y (nx5179), .A0 (nx5181), .A1 (nx5229), .S0 (nx5231)) ;
    mux21_ni ix5182 (.Y (nx5181), .A0 (nx5183), .A1 (nx5223), .S0 (nx5225)) ;
    mux21_ni ix5184 (.Y (nx5183), .A0 (nx5185), .A1 (nx5217), .S0 (nx5219)) ;
    mux21_ni ix5186 (.Y (nx5185), .A0 (nx5187), .A1 (nx5211), .S0 (nx5213)) ;
    mux21_ni ix5188 (.Y (nx5187), .A0 (nx5189), .A1 (nx5205), .S0 (nx5207)) ;
    mux21_ni ix5190 (.Y (nx5189), .A0 (nx5191), .A1 (nx5193), .S0 (nx2956)) ;
    nand02_2x ix5192 (.Y (nx5191), .A0 (input_b[1]), .A1 (input_a[2])) ;
    xnor2 ix2957 (.Y (nx2956), .A0 (nx2954), .A1 (nx5191)) ;
    inv02 ix5202 (.Y (nx5201), .A (input_b[2])) ;
    aoi22 ix5204 (.Y (nx5203), .A0 (input_b[3]), .A1 (input_a[0]), .B0 (
          input_b[2]), .B1 (input_a[1])) ;
    nand02_2x ix5206 (.Y (nx5205), .A0 (input_b[1]), .A1 (input_a[3])) ;
    xnor2 ix5208 (.Y (nx5207), .A0 (nx5209), .A1 (nx5205)) ;
    nand02_2x ix5212 (.Y (nx5211), .A0 (input_b[1]), .A1 (input_a[4])) ;
    xnor2 ix5214 (.Y (nx5213), .A0 (nx5215), .A1 (nx5211)) ;
    xnor2 ix5216 (.Y (nx5215), .A0 (nx4833), .A1 (nx4853)) ;
    nand02_2x ix5218 (.Y (nx5217), .A0 (input_b[1]), .A1 (input_a[5])) ;
    xnor2 ix5220 (.Y (nx5219), .A0 (nx5221), .A1 (nx5217)) ;
    xnor2 ix5222 (.Y (nx5221), .A0 (nx4831), .A1 (nx4869)) ;
    nand02_2x ix5224 (.Y (nx5223), .A0 (input_b[1]), .A1 (input_a[6])) ;
    xnor2 ix5226 (.Y (nx5225), .A0 (nx5227), .A1 (nx5223)) ;
    xnor2 ix5228 (.Y (nx5227), .A0 (nx4829), .A1 (nx4885)) ;
    nand02_2x ix5230 (.Y (nx5229), .A0 (input_b[1]), .A1 (input_a[7])) ;
    xnor2 ix5232 (.Y (nx5231), .A0 (nx5233), .A1 (nx5229)) ;
    xnor2 ix5234 (.Y (nx5233), .A0 (nx4827), .A1 (nx4899)) ;
    nand02_2x ix5236 (.Y (nx5235), .A0 (input_b[1]), .A1 (input_a[8])) ;
    xnor2 ix5238 (.Y (nx5237), .A0 (nx5239), .A1 (nx5235)) ;
    xnor2 ix5240 (.Y (nx5239), .A0 (nx4825), .A1 (nx4913)) ;
    nand02_2x ix5242 (.Y (nx5241), .A0 (input_b[1]), .A1 (input_a[9])) ;
    xnor2 ix5244 (.Y (nx5243), .A0 (nx5245), .A1 (nx5241)) ;
    xnor2 ix5246 (.Y (nx5245), .A0 (nx4823), .A1 (nx4927)) ;
    nand02_2x ix5248 (.Y (nx5247), .A0 (input_b[1]), .A1 (input_a[10])) ;
    xnor2 ix5250 (.Y (nx5249), .A0 (nx5251), .A1 (nx5247)) ;
    xnor2 ix5252 (.Y (nx5251), .A0 (nx4821), .A1 (nx4941)) ;
    nand02_2x ix5254 (.Y (nx5253), .A0 (input_b[1]), .A1 (input_a[11])) ;
    xnor2 ix5256 (.Y (nx5255), .A0 (nx5257), .A1 (nx5253)) ;
    xnor2 ix5258 (.Y (nx5257), .A0 (nx4819), .A1 (nx4955)) ;
    nand02_2x ix5260 (.Y (nx5259), .A0 (input_b[1]), .A1 (input_a[12])) ;
    xnor2 ix5262 (.Y (nx5261), .A0 (nx5263), .A1 (nx5259)) ;
    xnor2 ix5264 (.Y (nx5263), .A0 (nx4817), .A1 (nx4969)) ;
    nand02_2x ix5266 (.Y (nx5265), .A0 (input_b[1]), .A1 (input_a[13])) ;
    xnor2 ix5268 (.Y (nx5267), .A0 (nx5269), .A1 (nx5265)) ;
    xnor2 ix5270 (.Y (nx5269), .A0 (nx4815), .A1 (nx4983)) ;
    nand02_2x ix5272 (.Y (nx5271), .A0 (input_b[1]), .A1 (input_a[14])) ;
    xnor2 ix5274 (.Y (nx5273), .A0 (nx5275), .A1 (nx5271)) ;
    xnor2 ix5276 (.Y (nx5275), .A0 (nx4813), .A1 (nx4997)) ;
    nand02_2x ix5278 (.Y (nx5277), .A0 (input_b[1]), .A1 (input_a[15])) ;
    xnor2 ix5280 (.Y (nx5279), .A0 (nx5281), .A1 (nx5277)) ;
    xnor2 ix5282 (.Y (nx5281), .A0 (nx4811), .A1 (nx5011)) ;
    nand02_2x ix5284 (.Y (nx5283), .A0 (input_b[1]), .A1 (input_a[16])) ;
    xnor2 ix5286 (.Y (nx5285), .A0 (nx5287), .A1 (nx5283)) ;
    xnor2 ix5288 (.Y (nx5287), .A0 (nx4809), .A1 (nx5025)) ;
    nand02_2x ix5290 (.Y (nx5289), .A0 (input_b[1]), .A1 (input_a[17])) ;
    xnor2 ix5292 (.Y (nx5291), .A0 (nx5293), .A1 (nx5289)) ;
    xnor2 ix5294 (.Y (nx5293), .A0 (nx4807), .A1 (nx5039)) ;
    nand02_2x ix5296 (.Y (nx5295), .A0 (input_b[1]), .A1 (input_a[18])) ;
    xnor2 ix5298 (.Y (nx5297), .A0 (nx5299), .A1 (nx5295)) ;
    xnor2 ix5300 (.Y (nx5299), .A0 (nx4805), .A1 (nx5053)) ;
    nand02_2x ix5302 (.Y (nx5301), .A0 (input_b[1]), .A1 (input_a[19])) ;
    xnor2 ix5304 (.Y (nx5303), .A0 (nx5305), .A1 (nx5301)) ;
    xnor2 ix5306 (.Y (nx5305), .A0 (nx4803), .A1 (nx5067)) ;
    nand02_2x ix5308 (.Y (nx5307), .A0 (input_b[1]), .A1 (input_a[20])) ;
    xnor2 ix5310 (.Y (nx5309), .A0 (nx5311), .A1 (nx5307)) ;
    xnor2 ix5312 (.Y (nx5311), .A0 (nx4801), .A1 (nx5081)) ;
    xnor2 ix3321 (.Y (nx3320), .A0 (nx3316), .A1 (nx5151)) ;
    xnor2 ix3317 (.Y (nx3316), .A0 (nx4799), .A1 (nx3314)) ;
    xnor2 ix3919 (.Y (nx3918), .A0 (nx3914), .A1 (nx5321)) ;
    xnor2 ix3915 (.Y (nx3914), .A0 (nx4795), .A1 (nx3912)) ;
    nand02_2x ix5322 (.Y (nx5321), .A0 (input_b[1]), .A1 (input_a[22])) ;
    inv02 ix5324 (.Y (nx5323), .A (input_b[0])) ;
    mux21_ni ix5326 (.Y (nx5325), .A0 (nx5327), .A1 (nx5329), .S0 (nx3324)) ;
    nand02_2x ix5328 (.Y (nx5327), .A0 (input_b[0]), .A1 (input_a[22])) ;
    mux21_ni ix5330 (.Y (nx5329), .A0 (nx5331), .A1 (nx5491), .S0 (nx5493)) ;
    mux21_ni ix5332 (.Y (nx5331), .A0 (nx5333), .A1 (nx5485), .S0 (nx5487)) ;
    mux21_ni ix5334 (.Y (nx5333), .A0 (nx5335), .A1 (nx5479), .S0 (nx5481)) ;
    mux21_ni ix5336 (.Y (nx5335), .A0 (nx5337), .A1 (nx5473), .S0 (nx5475)) ;
    mux21_ni ix5338 (.Y (nx5337), .A0 (nx5339), .A1 (nx5467), .S0 (nx5469)) ;
    mux21_ni ix5340 (.Y (nx5339), .A0 (nx5341), .A1 (nx5461), .S0 (nx5463)) ;
    mux21_ni ix5342 (.Y (nx5341), .A0 (nx5343), .A1 (nx5455), .S0 (nx5457)) ;
    mux21_ni ix5344 (.Y (nx5343), .A0 (nx5345), .A1 (nx5449), .S0 (nx5451)) ;
    mux21_ni ix5346 (.Y (nx5345), .A0 (nx5347), .A1 (nx5443), .S0 (nx5445)) ;
    mux21_ni ix5348 (.Y (nx5347), .A0 (nx5349), .A1 (nx5437), .S0 (nx5439)) ;
    mux21_ni ix5350 (.Y (nx5349), .A0 (nx5351), .A1 (nx5431), .S0 (nx5433)) ;
    mux21_ni ix5352 (.Y (nx5351), .A0 (nx5353), .A1 (nx5425), .S0 (nx5427)) ;
    mux21_ni ix5354 (.Y (nx5353), .A0 (nx5355), .A1 (nx5419), .S0 (nx5421)) ;
    mux21_ni ix5356 (.Y (nx5355), .A0 (nx5357), .A1 (nx5413), .S0 (nx5415)) ;
    mux21_ni ix5358 (.Y (nx5357), .A0 (nx5359), .A1 (nx5407), .S0 (nx5409)) ;
    mux21_ni ix5360 (.Y (nx5359), .A0 (nx5361), .A1 (nx5401), .S0 (nx5403)) ;
    mux21_ni ix5362 (.Y (nx5361), .A0 (nx5363), .A1 (nx5395), .S0 (nx5397)) ;
    mux21_ni ix5364 (.Y (nx5363), .A0 (nx5365), .A1 (nx5389), .S0 (nx5391)) ;
    mux21_ni ix5366 (.Y (nx5365), .A0 (nx5367), .A1 (nx5383), .S0 (nx5385)) ;
    mux21_ni ix5368 (.Y (nx5367), .A0 (nx5369), .A1 (nx5371), .S0 (nx3532)) ;
    nand02_2x ix5370 (.Y (nx5369), .A0 (input_b[0]), .A1 (input_a[2])) ;
    xnor2 ix3533 (.Y (nx3532), .A0 (nx3530), .A1 (nx5369)) ;
    inv02 ix5380 (.Y (nx5379), .A (input_b[1])) ;
    aoi22 ix5382 (.Y (nx5381), .A0 (input_b[2]), .A1 (input_a[0]), .B0 (
          input_b[1]), .B1 (input_a[1])) ;
    nand02_2x ix5384 (.Y (nx5383), .A0 (input_b[0]), .A1 (input_a[3])) ;
    xnor2 ix5386 (.Y (nx5385), .A0 (nx5387), .A1 (nx5383)) ;
    nand02_2x ix5390 (.Y (nx5389), .A0 (input_b[0]), .A1 (input_a[4])) ;
    xnor2 ix5392 (.Y (nx5391), .A0 (nx5393), .A1 (nx5389)) ;
    xnor2 ix5394 (.Y (nx5393), .A0 (nx5189), .A1 (nx5207)) ;
    nand02_2x ix5396 (.Y (nx5395), .A0 (input_b[0]), .A1 (input_a[5])) ;
    xnor2 ix5398 (.Y (nx5397), .A0 (nx5399), .A1 (nx5395)) ;
    xnor2 ix5400 (.Y (nx5399), .A0 (nx5187), .A1 (nx5213)) ;
    nand02_2x ix5402 (.Y (nx5401), .A0 (input_b[0]), .A1 (input_a[6])) ;
    xnor2 ix5404 (.Y (nx5403), .A0 (nx5405), .A1 (nx5401)) ;
    xnor2 ix5406 (.Y (nx5405), .A0 (nx5185), .A1 (nx5219)) ;
    nand02_2x ix5408 (.Y (nx5407), .A0 (input_b[0]), .A1 (input_a[7])) ;
    xnor2 ix5410 (.Y (nx5409), .A0 (nx5411), .A1 (nx5407)) ;
    xnor2 ix5412 (.Y (nx5411), .A0 (nx5183), .A1 (nx5225)) ;
    nand02_2x ix5414 (.Y (nx5413), .A0 (input_b[0]), .A1 (input_a[8])) ;
    xnor2 ix5416 (.Y (nx5415), .A0 (nx5417), .A1 (nx5413)) ;
    xnor2 ix5418 (.Y (nx5417), .A0 (nx5181), .A1 (nx5231)) ;
    nand02_2x ix5420 (.Y (nx5419), .A0 (input_b[0]), .A1 (input_a[9])) ;
    xnor2 ix5422 (.Y (nx5421), .A0 (nx5423), .A1 (nx5419)) ;
    xnor2 ix5424 (.Y (nx5423), .A0 (nx5179), .A1 (nx5237)) ;
    nand02_2x ix5426 (.Y (nx5425), .A0 (input_b[0]), .A1 (input_a[10])) ;
    xnor2 ix5428 (.Y (nx5427), .A0 (nx5429), .A1 (nx5425)) ;
    xnor2 ix5430 (.Y (nx5429), .A0 (nx5177), .A1 (nx5243)) ;
    nand02_2x ix5432 (.Y (nx5431), .A0 (input_b[0]), .A1 (input_a[11])) ;
    xnor2 ix5434 (.Y (nx5433), .A0 (nx5435), .A1 (nx5431)) ;
    xnor2 ix5436 (.Y (nx5435), .A0 (nx5175), .A1 (nx5249)) ;
    nand02_2x ix5438 (.Y (nx5437), .A0 (input_b[0]), .A1 (input_a[12])) ;
    xnor2 ix5440 (.Y (nx5439), .A0 (nx5441), .A1 (nx5437)) ;
    xnor2 ix5442 (.Y (nx5441), .A0 (nx5173), .A1 (nx5255)) ;
    nand02_2x ix5444 (.Y (nx5443), .A0 (input_b[0]), .A1 (input_a[13])) ;
    xnor2 ix5446 (.Y (nx5445), .A0 (nx5447), .A1 (nx5443)) ;
    xnor2 ix5448 (.Y (nx5447), .A0 (nx5171), .A1 (nx5261)) ;
    nand02_2x ix5450 (.Y (nx5449), .A0 (input_b[0]), .A1 (input_a[14])) ;
    xnor2 ix5452 (.Y (nx5451), .A0 (nx5453), .A1 (nx5449)) ;
    xnor2 ix5454 (.Y (nx5453), .A0 (nx5169), .A1 (nx5267)) ;
    nand02_2x ix5456 (.Y (nx5455), .A0 (input_b[0]), .A1 (input_a[15])) ;
    xnor2 ix5458 (.Y (nx5457), .A0 (nx5459), .A1 (nx5455)) ;
    xnor2 ix5460 (.Y (nx5459), .A0 (nx5167), .A1 (nx5273)) ;
    nand02_2x ix5462 (.Y (nx5461), .A0 (input_b[0]), .A1 (input_a[16])) ;
    xnor2 ix5464 (.Y (nx5463), .A0 (nx5465), .A1 (nx5461)) ;
    xnor2 ix5466 (.Y (nx5465), .A0 (nx5165), .A1 (nx5279)) ;
    nand02_2x ix5468 (.Y (nx5467), .A0 (input_b[0]), .A1 (input_a[17])) ;
    xnor2 ix5470 (.Y (nx5469), .A0 (nx5471), .A1 (nx5467)) ;
    xnor2 ix5472 (.Y (nx5471), .A0 (nx5163), .A1 (nx5285)) ;
    nand02_2x ix5474 (.Y (nx5473), .A0 (input_b[0]), .A1 (input_a[18])) ;
    xnor2 ix5476 (.Y (nx5475), .A0 (nx5477), .A1 (nx5473)) ;
    xnor2 ix5478 (.Y (nx5477), .A0 (nx5161), .A1 (nx5291)) ;
    nand02_2x ix5480 (.Y (nx5479), .A0 (input_b[0]), .A1 (input_a[19])) ;
    xnor2 ix5482 (.Y (nx5481), .A0 (nx5483), .A1 (nx5479)) ;
    xnor2 ix5484 (.Y (nx5483), .A0 (nx5159), .A1 (nx5297)) ;
    nand02_2x ix5486 (.Y (nx5485), .A0 (input_b[0]), .A1 (input_a[20])) ;
    xnor2 ix5488 (.Y (nx5487), .A0 (nx5489), .A1 (nx5485)) ;
    xnor2 ix5490 (.Y (nx5489), .A0 (nx5157), .A1 (nx5303)) ;
    nand02_2x ix5492 (.Y (nx5491), .A0 (input_b[0]), .A1 (input_a[21])) ;
    xnor2 ix5494 (.Y (nx5493), .A0 (nx5495), .A1 (nx5491)) ;
    xnor2 ix5496 (.Y (nx5495), .A0 (nx5155), .A1 (nx5309)) ;
    xnor2 ix3325 (.Y (nx3324), .A0 (nx3322), .A1 (nx5327)) ;
    xnor2 ix3323 (.Y (nx3322), .A0 (nx5153), .A1 (nx3320)) ;
    xnor2 ix5502 (.Y (nx5501), .A0 (input_b[0]), .A1 (nx3920)) ;
    xnor2 ix3921 (.Y (nx3920), .A0 (nx5149), .A1 (nx3918)) ;
    xnor2 ix7827 (.Y (nx7826), .A0 (nx5507), .A1 (nx7794)) ;
    mux21_ni ix5508 (.Y (nx5507), .A0 (nx5321), .A1 (nx5149), .S0 (nx3918)) ;
    xnor2 ix7795 (.Y (nx7794), .A0 (input_b[1]), .A1 (nx5511)) ;
    xnor2 ix5512 (.Y (nx5511), .A0 (nx4791), .A1 (nx5119)) ;
    xnor2 ix7813 (.Y (nx7812), .A0 (nx7810), .A1 (nx4787)) ;
    oai22 ix7811 (.Y (nx7810), .A0 (nx5507), .A1 (nx5517), .B0 (nx5511), .B1 (
          nx5379)) ;
    xnor2 ix7749 (.Y (nx7748), .A0 (nx5521), .A1 (nx7696)) ;
    mux21_ni ix5522 (.Y (nx5521), .A0 (nx5141), .A1 (nx5135), .S0 (nx7706)) ;
    xnor2 ix7697 (.Y (nx7696), .A0 (input_b[3]), .A1 (nx5525)) ;
    xnor2 ix5526 (.Y (nx5525), .A0 (nx4431), .A1 (nx4759)) ;
    xnor2 ix5528 (.Y (nx5527), .A0 (nx7782), .A1 (nx7748)) ;
    oai22 ix7783 (.Y (nx7782), .A0 (nx5531), .A1 (nx5201), .B0 (nx4789), .B1 (
          nx5131)) ;
    xnor2 ix7743 (.Y (nx7742), .A0 (nx7740), .A1 (nx5539)) ;
    oai22 ix7741 (.Y (nx7740), .A0 (nx5521), .A1 (nx5537), .B0 (nx5525), .B1 (
          nx4845)) ;
    xnor2 ix5540 (.Y (nx5539), .A0 (nx4429), .A1 (nx4771)) ;
    xnor2 ix7623 (.Y (nx7622), .A0 (nx5543), .A1 (nx7542)) ;
    mux21_ni ix5544 (.Y (nx5543), .A0 (nx4781), .A1 (nx4775), .S0 (nx7552)) ;
    xnor2 ix7543 (.Y (nx7542), .A0 (input_b[5]), .A1 (nx5547)) ;
    xnor2 ix5548 (.Y (nx5547), .A0 (nx4071), .A1 (nx4399)) ;
    xnor2 ix5550 (.Y (nx5549), .A0 (nx7684), .A1 (nx7622)) ;
    oai22 ix7685 (.Y (nx7684), .A0 (nx5553), .A1 (nx4847), .B0 (nx4429), .B1 (
          nx4771)) ;
    xnor2 ix7617 (.Y (nx7616), .A0 (nx7614), .A1 (nx4067)) ;
    oai22 ix7615 (.Y (nx7614), .A0 (nx5543), .A1 (nx5559), .B0 (nx5547), .B1 (
          nx4487)) ;
    mux21_ni ix5564 (.Y (nx5563), .A0 (nx4421), .A1 (nx4415), .S0 (nx7342)) ;
    xnor2 ix7333 (.Y (nx7332), .A0 (input_b[7]), .A1 (nx5567)) ;
    xnor2 ix5568 (.Y (nx5567), .A0 (nx3711), .A1 (nx4039)) ;
    xnor2 ix5570 (.Y (nx5569), .A0 (nx7530), .A1 (nx7440)) ;
    oai22 ix7531 (.Y (nx7530), .A0 (nx5573), .A1 (nx4489), .B0 (nx4069), .B1 (
          nx4411)) ;
    xnor2 ix7441 (.Y (nx7440), .A0 (nx5563), .A1 (nx7332)) ;
    xnor2 ix7435 (.Y (nx7434), .A0 (nx7432), .A1 (nx3707)) ;
    oai22 ix7433 (.Y (nx7432), .A0 (nx5563), .A1 (nx5581), .B0 (nx5567), .B1 (
          nx4129)) ;
    xnor2 ix7203 (.Y (nx7202), .A0 (nx5585), .A1 (nx7066)) ;
    mux21_ni ix5586 (.Y (nx5585), .A0 (nx4061), .A1 (nx4055), .S0 (nx7076)) ;
    xnor2 ix7067 (.Y (nx7066), .A0 (input_b[9]), .A1 (nx5589)) ;
    xnor2 ix5590 (.Y (nx5589), .A0 (nx3351), .A1 (nx3679)) ;
    xnor2 ix5592 (.Y (nx5591), .A0 (nx7320), .A1 (nx7202)) ;
    oai22 ix7321 (.Y (nx7320), .A0 (nx5595), .A1 (nx4131), .B0 (nx3709), .B1 (
          nx4051)) ;
    xnor2 ix7197 (.Y (nx7196), .A0 (nx7194), .A1 (nx5603)) ;
    oai22 ix7195 (.Y (nx7194), .A0 (nx5585), .A1 (nx5601), .B0 (nx5589), .B1 (
          nx3771)) ;
    xnor2 ix5604 (.Y (nx5603), .A0 (nx3349), .A1 (nx3691)) ;
    xnor2 ix6909 (.Y (nx6908), .A0 (nx5607), .A1 (nx6744)) ;
    mux21_ni ix5608 (.Y (nx5607), .A0 (nx3701), .A1 (nx3695), .S0 (nx6754)) ;
    xnor2 ix6745 (.Y (nx6744), .A0 (input_b[11]), .A1 (nx5611)) ;
    xnor2 ix5612 (.Y (nx5611), .A0 (nx2991), .A1 (nx3319)) ;
    xnor2 ix5614 (.Y (nx5613), .A0 (nx7054), .A1 (nx6908)) ;
    oai22 ix7055 (.Y (nx7054), .A0 (nx3349), .A1 (nx3691), .B0 (nx5617), .B1 (
          nx3773)) ;
    xnor2 ix6903 (.Y (nx6902), .A0 (nx6900), .A1 (nx2987)) ;
    oai22 ix6901 (.Y (nx6900), .A0 (nx5607), .A1 (nx5623), .B0 (nx5611), .B1 (
          nx3413)) ;
    mux21_ni ix5628 (.Y (nx5627), .A0 (nx3341), .A1 (nx3335), .S0 (nx6376)) ;
    xnor2 ix6367 (.Y (nx6366), .A0 (input_b[13]), .A1 (nx5631)) ;
    xnor2 ix5632 (.Y (nx5631), .A0 (nx2631), .A1 (nx2959)) ;
    xnor2 ix5634 (.Y (nx5633), .A0 (nx6732), .A1 (nx6558)) ;
    oai22 ix6733 (.Y (nx6732), .A0 (nx2989), .A1 (nx3331), .B0 (nx5637), .B1 (
          nx3415)) ;
    xnor2 ix6559 (.Y (nx6558), .A0 (nx5627), .A1 (nx6366)) ;
    xnor2 ix6553 (.Y (nx6552), .A0 (nx6550), .A1 (nx2627)) ;
    oai22 ix6551 (.Y (nx6550), .A0 (nx5627), .A1 (nx5645), .B0 (nx5631), .B1 (
          nx3055)) ;
    xnor2 ix6153 (.Y (nx6152), .A0 (nx5649), .A1 (nx5932)) ;
    mux21_ni ix5650 (.Y (nx5649), .A0 (nx2981), .A1 (nx2975), .S0 (nx5942)) ;
    xnor2 ix5933 (.Y (nx5932), .A0 (input_b[15]), .A1 (nx5653)) ;
    xnor2 ix5654 (.Y (nx5653), .A0 (nx2271), .A1 (nx2599)) ;
    xnor2 ix5656 (.Y (nx5655), .A0 (nx6354), .A1 (nx6152)) ;
    oai22 ix6355 (.Y (nx6354), .A0 (nx2629), .A1 (nx2971), .B0 (nx5659), .B1 (
          nx3057)) ;
    xnor2 ix6147 (.Y (nx6146), .A0 (nx6144), .A1 (nx5667)) ;
    oai22 ix6145 (.Y (nx6144), .A0 (nx5649), .A1 (nx5665), .B0 (nx5653), .B1 (
          nx2697)) ;
    xnor2 ix5668 (.Y (nx5667), .A0 (nx2269), .A1 (nx2611)) ;
    xnor2 ix5691 (.Y (nx5690), .A0 (nx5671), .A1 (nx5442)) ;
    mux21_ni ix5672 (.Y (nx5671), .A0 (nx2621), .A1 (nx2615), .S0 (nx5452)) ;
    xnor2 ix5443 (.Y (nx5442), .A0 (input_b[17]), .A1 (nx5675)) ;
    xnor2 ix5676 (.Y (nx5675), .A0 (nx1911), .A1 (nx2239)) ;
    xnor2 ix5678 (.Y (nx5677), .A0 (nx5920), .A1 (nx5690)) ;
    oai22 ix5921 (.Y (nx5920), .A0 (nx2269), .A1 (nx2611), .B0 (nx5681), .B1 (
          nx2699)) ;
    xnor2 ix5685 (.Y (nx5684), .A0 (nx5682), .A1 (nx1907)) ;
    oai22 ix5683 (.Y (nx5682), .A0 (nx5671), .A1 (nx5687), .B0 (nx5675), .B1 (
          nx2339)) ;
    mux21_ni ix5692 (.Y (nx5691), .A0 (nx2261), .A1 (nx2255), .S0 (nx4906)) ;
    xnor2 ix4897 (.Y (nx4896), .A0 (input_b[19]), .A1 (nx5695)) ;
    xnor2 ix5696 (.Y (nx5695), .A0 (nx1529), .A1 (nx1877)) ;
    xnor2 ix5698 (.Y (nx5697), .A0 (nx5430), .A1 (nx5172)) ;
    oai22 ix5431 (.Y (nx5430), .A0 (nx1909), .A1 (nx2251), .B0 (nx5701), .B1 (
          nx2341)) ;
    xnor2 ix5173 (.Y (nx5172), .A0 (nx5691), .A1 (nx4896)) ;
    xnor2 ix5167 (.Y (nx5166), .A0 (nx5164), .A1 (nx1525)) ;
    oai22 ix5165 (.Y (nx5164), .A0 (nx5691), .A1 (nx5709), .B0 (nx5695), .B1 (
          nx1981)) ;
    xnor2 ix4599 (.Y (nx4598), .A0 (nx5713), .A1 (nx4294)) ;
    mux21_ni ix5714 (.Y (nx5713), .A0 (nx1901), .A1 (nx1893), .S0 (nx4304)) ;
    xnor2 ix4295 (.Y (nx4294), .A0 (input_b[21]), .A1 (nx5717)) ;
    xnor2 ix5718 (.Y (nx5717), .A0 (nx6389), .A1 (nx4030)) ;
    xnor2 ix5720 (.Y (nx5719), .A0 (nx4884), .A1 (nx4598)) ;
    oai22 ix4885 (.Y (nx4884), .A0 (nx1527), .A1 (nx1889), .B0 (nx5723), .B1 (
          nx1983)) ;
    xnor2 ix4593 (.Y (nx4592), .A0 (nx4590), .A1 (nx5731)) ;
    oai22 ix4591 (.Y (nx4590), .A0 (nx5713), .A1 (nx5729), .B0 (nx5717), .B1 (
          nx1609)) ;
    xnor2 ix5732 (.Y (nx5731), .A0 (nx1349), .A1 (nx1519)) ;
    oai21 ix4289 (.Y (nx4288), .A0 (nx1349), .A1 (nx1519), .B0 (nx1517)) ;
    nand02_2x ix5736 (.Y (nx5735), .A0 (nx7920), .A1 (nx8012)) ;
    xnor2 ix7921 (.Y (nx7920), .A0 (nx4288), .A1 (nx7912)) ;
    nor02ii ix8013 (.Y (nx8012), .A0 (nx5741), .A1 (nx8010)) ;
    xnor2 ix5742 (.Y (nx5741), .A0 (nx7908), .A1 (nx4592)) ;
    nor02_2x ix8011 (.Y (nx8010), .A0 (nx5745), .A1 (nx5749)) ;
    xnor2 ix5746 (.Y (nx5745), .A0 (nx5747), .A1 (nx5719)) ;
    mux21_ni ix5748 (.Y (nx5747), .A0 (nx1525), .A1 (nx1903), .S0 (nx5166)) ;
    nand02_2x ix5750 (.Y (nx5749), .A0 (nx7926), .A1 (nx6403)) ;
    xnor2 ix7927 (.Y (nx7926), .A0 (nx1903), .A1 (nx5166)) ;
    nor02ii ix8007 (.Y (nx8006), .A0 (nx5755), .A1 (nx8004)) ;
    xnor2 ix5756 (.Y (nx5755), .A0 (nx1905), .A1 (nx5697)) ;
    nor02_2x ix8005 (.Y (nx8004), .A0 (nx5759), .A1 (nx5763)) ;
    xnor2 ix5760 (.Y (nx5759), .A0 (nx7892), .A1 (nx5684)) ;
    mux21_ni ix7893 (.Y (nx7892), .A0 (nx7888), .A1 (nx5690), .S0 (nx5677)) ;
    nand02_2x ix5764 (.Y (nx5763), .A0 (nx7932), .A1 (nx6401)) ;
    xnor2 ix7933 (.Y (nx7932), .A0 (nx7888), .A1 (nx5677)) ;
    nor02ii ix8001 (.Y (nx8000), .A0 (nx5769), .A1 (nx7998)) ;
    xnor2 ix5770 (.Y (nx5769), .A0 (nx7884), .A1 (nx6146)) ;
    nor02_2x ix7999 (.Y (nx7998), .A0 (nx5773), .A1 (nx5777)) ;
    xnor2 ix5774 (.Y (nx5773), .A0 (nx5775), .A1 (nx5655)) ;
    mux21_ni ix5776 (.Y (nx5775), .A0 (nx2627), .A1 (nx2983), .S0 (nx6552)) ;
    nand02_2x ix5778 (.Y (nx5777), .A0 (nx7938), .A1 (nx6399)) ;
    xnor2 ix7939 (.Y (nx7938), .A0 (nx2983), .A1 (nx6552)) ;
    nor02ii ix7995 (.Y (nx7994), .A0 (nx5783), .A1 (nx7992)) ;
    xnor2 ix5784 (.Y (nx5783), .A0 (nx2985), .A1 (nx5633)) ;
    nor02_2x ix7993 (.Y (nx7992), .A0 (nx5787), .A1 (nx5791)) ;
    xnor2 ix5788 (.Y (nx5787), .A0 (nx7868), .A1 (nx6902)) ;
    mux21_ni ix7869 (.Y (nx7868), .A0 (nx7864), .A1 (nx6908), .S0 (nx5613)) ;
    nand02_2x ix5792 (.Y (nx5791), .A0 (nx7944), .A1 (nx6397)) ;
    xnor2 ix7945 (.Y (nx7944), .A0 (nx7864), .A1 (nx5613)) ;
    nor02ii ix7989 (.Y (nx7988), .A0 (nx5797), .A1 (nx7986)) ;
    xnor2 ix5798 (.Y (nx5797), .A0 (nx7860), .A1 (nx7196)) ;
    nor02_2x ix7987 (.Y (nx7986), .A0 (nx5801), .A1 (nx5805)) ;
    xnor2 ix5802 (.Y (nx5801), .A0 (nx5803), .A1 (nx5591)) ;
    mux21_ni ix5804 (.Y (nx5803), .A0 (nx3707), .A1 (nx4063), .S0 (nx7434)) ;
    nand02_2x ix5806 (.Y (nx5805), .A0 (nx7950), .A1 (nx6395)) ;
    xnor2 ix7951 (.Y (nx7950), .A0 (nx4063), .A1 (nx7434)) ;
    nor02ii ix7983 (.Y (nx7982), .A0 (nx5811), .A1 (nx7980)) ;
    xnor2 ix5812 (.Y (nx5811), .A0 (nx4065), .A1 (nx5569)) ;
    nor02_2x ix7981 (.Y (nx7980), .A0 (nx5815), .A1 (nx5819)) ;
    xnor2 ix5816 (.Y (nx5815), .A0 (nx7844), .A1 (nx7616)) ;
    mux21_ni ix7845 (.Y (nx7844), .A0 (nx7840), .A1 (nx7622), .S0 (nx5549)) ;
    nand02_2x ix5820 (.Y (nx5819), .A0 (nx7956), .A1 (nx6393)) ;
    xnor2 ix7957 (.Y (nx7956), .A0 (nx7840), .A1 (nx5549)) ;
    nor02ii ix7977 (.Y (nx7976), .A0 (nx5825), .A1 (nx7974)) ;
    xnor2 ix5826 (.Y (nx5825), .A0 (nx7836), .A1 (nx7742)) ;
    nor02_2x ix7975 (.Y (nx7974), .A0 (nx5829), .A1 (nx5833)) ;
    xnor2 ix5830 (.Y (nx5829), .A0 (nx5831), .A1 (nx5527)) ;
    mux21_ni ix5832 (.Y (nx5831), .A0 (nx4787), .A1 (nx5143), .S0 (nx7812)) ;
    nand02_2x ix5834 (.Y (nx5833), .A0 (nx7962), .A1 (nx6391)) ;
    xnor2 ix7963 (.Y (nx7962), .A0 (nx5143), .A1 (nx7812)) ;
    nor02ii ix7971 (.Y (nx7970), .A0 (nx5839), .A1 (nx4020)) ;
    xnor2 ix5840 (.Y (nx5839), .A0 (nx7824), .A1 (nx7826)) ;
    nor02_2x ix4021 (.Y (nx4020), .A0 (nx5843), .A1 (nx5845)) ;
    xnor2 ix5844 (.Y (nx5843), .A0 (nx5325), .A1 (nx5501)) ;
    nand04 ix5846 (.Y (nx5845), .A0 (nx3946), .A1 (nx3968), .A2 (nx3992), .A3 (
           nx4014)) ;
    nor04 ix3947 (.Y (nx3946), .A0 (nx5849), .A1 (nx5853), .A2 (nx5855), .A3 (
          nx5857)) ;
    nand04 ix5850 (.Y (nx5849), .A0 (input_b[0]), .A1 (input_a[0]), .A2 (nx5371)
           , .A3 (nx3928)) ;
    xnor2 ix3929 (.Y (nx3928), .A0 (nx5329), .A1 (nx3324)) ;
    xnor2 ix5854 (.Y (nx5853), .A0 (nx5335), .A1 (nx5481)) ;
    xnor2 ix5856 (.Y (nx5855), .A0 (nx5331), .A1 (nx5493)) ;
    xnor2 ix5858 (.Y (nx5857), .A0 (nx5333), .A1 (nx5487)) ;
    nor04 ix3969 (.Y (nx3968), .A0 (nx5861), .A1 (nx5863), .A2 (nx5865), .A3 (
          nx5867)) ;
    xnor2 ix5862 (.Y (nx5861), .A0 (nx5341), .A1 (nx5463)) ;
    xnor2 ix5864 (.Y (nx5863), .A0 (nx5337), .A1 (nx5475)) ;
    xnor2 ix5866 (.Y (nx5865), .A0 (nx5339), .A1 (nx5469)) ;
    or03 ix5868 (.Y (nx5867), .A0 (nx5869), .A1 (nx5871), .A2 (nx5873)) ;
    xnor2 ix5870 (.Y (nx5869), .A0 (nx5347), .A1 (nx5445)) ;
    xnor2 ix5872 (.Y (nx5871), .A0 (nx5343), .A1 (nx5457)) ;
    xnor2 ix5874 (.Y (nx5873), .A0 (nx5345), .A1 (nx5451)) ;
    nor04 ix3993 (.Y (nx3992), .A0 (nx5877), .A1 (nx5879), .A2 (nx5881), .A3 (
          nx5883)) ;
    xnor2 ix5878 (.Y (nx5877), .A0 (nx5353), .A1 (nx5427)) ;
    xnor2 ix5880 (.Y (nx5879), .A0 (nx5349), .A1 (nx5439)) ;
    xnor2 ix5882 (.Y (nx5881), .A0 (nx5351), .A1 (nx5433)) ;
    or03 ix5884 (.Y (nx5883), .A0 (nx5885), .A1 (nx5887), .A2 (nx5889)) ;
    xnor2 ix5886 (.Y (nx5885), .A0 (nx5359), .A1 (nx5409)) ;
    xnor2 ix5888 (.Y (nx5887), .A0 (nx5355), .A1 (nx5421)) ;
    xnor2 ix5890 (.Y (nx5889), .A0 (nx5357), .A1 (nx5415)) ;
    nor04 ix4015 (.Y (nx4014), .A0 (nx5893), .A1 (nx5895), .A2 (nx5897), .A3 (
          nx5899)) ;
    xnor2 ix5894 (.Y (nx5893), .A0 (nx5365), .A1 (nx5391)) ;
    xnor2 ix5896 (.Y (nx5895), .A0 (nx5361), .A1 (nx5403)) ;
    xnor2 ix5898 (.Y (nx5897), .A0 (nx5363), .A1 (nx5397)) ;
    oai21 ix5900 (.Y (nx5899), .A0 (input_a[1]), .A1 (input_b[1]), .B0 (nx4010)
          ) ;
    nor02_2x ix4011 (.Y (nx4010), .A0 (nx5903), .A1 (nx5905)) ;
    xnor2 ix5904 (.Y (nx5903), .A0 (nx5367), .A1 (nx5385)) ;
    xnor2 ix8733 (.Y (nx8732), .A0 (nx6427), .A1 (nx1293)) ;
    xnor2 ix8721 (.Y (nx8720), .A0 (nx8666), .A1 (nx1285)) ;
    nor03 ix8773 (.Y (underflow), .A0 (nx1245), .A1 (input_a[30]), .A2 (
          input_b[30])) ;
    oai22 ix253 (.Y (nx252), .A0 (nx5919), .A1 (nx5929), .B0 (nx5939), .B1 (
          nx5949)) ;
    nand04 ix5920 (.Y (nx5919), .A0 (nx138), .A1 (nx152), .A2 (nx168), .A3 (
           nx182)) ;
    nor04 ix139 (.Y (nx138), .A0 (input_b[0]), .A1 (input_b[1]), .A2 (input_b[2]
          ), .A3 (input_b[3])) ;
    nor04 ix153 (.Y (nx152), .A0 (input_b[4]), .A1 (input_b[5]), .A2 (input_b[6]
          ), .A3 (input_b[7])) ;
    nor04 ix169 (.Y (nx168), .A0 (input_b[8]), .A1 (input_b[9]), .A2 (
          input_b[10]), .A3 (input_b[11])) ;
    nor04 ix183 (.Y (nx182), .A0 (input_b[12]), .A1 (input_b[13]), .A2 (
          input_b[14]), .A3 (input_b[15])) ;
    nand04 ix5930 (.Y (nx5929), .A0 (nx200), .A1 (nx214), .A2 (nx230), .A3 (
           nx244)) ;
    nor04 ix201 (.Y (nx200), .A0 (input_b[16]), .A1 (input_b[17]), .A2 (
          input_b[18]), .A3 (input_b[19])) ;
    nor04 ix215 (.Y (nx214), .A0 (input_b[20]), .A1 (input_b[21]), .A2 (
          input_b[22]), .A3 (input_b[23])) ;
    nor04 ix231 (.Y (nx230), .A0 (input_b[24]), .A1 (input_b[25]), .A2 (
          input_b[26]), .A3 (input_b[27])) ;
    nor04 ix245 (.Y (nx244), .A0 (input_b[28]), .A1 (input_b[29]), .A2 (
          input_b[30]), .A3 (input_b[31])) ;
    nand04 ix5940 (.Y (nx5939), .A0 (nx12), .A1 (nx26), .A2 (nx42), .A3 (nx56)
           ) ;
    nor04 ix13 (.Y (nx12), .A0 (input_a[0]), .A1 (input_a[1]), .A2 (input_a[2])
          , .A3 (input_a[3])) ;
    nor04 ix27 (.Y (nx26), .A0 (input_a[4]), .A1 (input_a[5]), .A2 (input_a[6])
          , .A3 (input_a[7])) ;
    nor04 ix43 (.Y (nx42), .A0 (input_a[8]), .A1 (input_a[9]), .A2 (input_a[10])
          , .A3 (input_a[11])) ;
    nor04 ix57 (.Y (nx56), .A0 (input_a[12]), .A1 (input_a[13]), .A2 (
          input_a[14]), .A3 (input_a[15])) ;
    nand04 ix5950 (.Y (nx5949), .A0 (nx74), .A1 (nx88), .A2 (nx104), .A3 (nx118)
           ) ;
    nor04 ix75 (.Y (nx74), .A0 (input_a[16]), .A1 (input_a[17]), .A2 (
          input_a[18]), .A3 (input_a[19])) ;
    nor04 ix89 (.Y (nx88), .A0 (input_a[20]), .A1 (input_a[21]), .A2 (
          input_a[22]), .A3 (input_a[23])) ;
    nor04 ix105 (.Y (nx104), .A0 (input_a[24]), .A1 (input_a[25]), .A2 (
          input_a[26]), .A3 (input_a[27])) ;
    nor04 ix119 (.Y (nx118), .A0 (input_a[28]), .A1 (input_a[29]), .A2 (
          input_a[30]), .A3 (input_a[31])) ;
    xnor2 ix8029 (.Y (nx8028), .A0 (nx5839), .A1 (nx4020)) ;
    xnor2 ix5964 (.Y (nx5963), .A0 (nx5843), .A1 (nx5845)) ;
    aoi21 ix5968 (.Y (nx5967), .A0 (nx6405), .A1 (nx8054), .B0 (nx8048)) ;
    nor03 ix8049 (.Y (nx8048), .A0 (nx5975), .A1 (nx6405), .A2 (nx8040)) ;
    nor02ii ix5976 (.Y (nx5975), .A0 (nx8028), .A1 (nx5963)) ;
    nor02ii ix8041 (.Y (nx8040), .A0 (nx5963), .A1 (nx8028)) ;
    aoi21 ix5982 (.Y (nx5981), .A0 (nx6405), .A1 (nx8080), .B0 (nx8074)) ;
    nor03 ix8075 (.Y (nx8074), .A0 (nx5987), .A1 (nx6405), .A2 (nx8066)) ;
    nor02ii ix5988 (.Y (nx5987), .A0 (nx8040), .A1 (nx5989)) ;
    xnor2 ix5990 (.Y (nx5989), .A0 (nx7962), .A1 (nx6391)) ;
    nor02ii ix8067 (.Y (nx8066), .A0 (nx5989), .A1 (nx8040)) ;
    aoi21 ix5996 (.Y (nx5995), .A0 (nx6405), .A1 (nx8106), .B0 (nx8100)) ;
    xnor2 ix8107 (.Y (nx8106), .A0 (nx5825), .A1 (nx7974)) ;
    nor03 ix8101 (.Y (nx8100), .A0 (nx6001), .A1 (nx6405), .A2 (nx6413)) ;
    nor02ii ix6002 (.Y (nx6001), .A0 (nx8066), .A1 (nx6003)) ;
    xnor2 ix6004 (.Y (nx6003), .A0 (nx5829), .A1 (nx5833)) ;
    nor02ii ix8093 (.Y (nx8092), .A0 (nx6003), .A1 (nx8066)) ;
    oai22 ix8137 (.Y (nx8136), .A0 (nx6433), .A1 (nx6011), .B0 (nx6013), .B1 (
          nx6015)) ;
    xnor2 ix6012 (.Y (nx6011), .A0 (nx7956), .A1 (nx6393)) ;
    nor02_2x ix6014 (.Y (nx6013), .A0 (nx6413), .A1 (nx8106)) ;
    nand02_2x ix6016 (.Y (nx6015), .A0 (nx6433), .A1 (nx6017)) ;
    nand02_2x ix6018 (.Y (nx6017), .A0 (nx8106), .A1 (nx6413)) ;
    aoi22 ix6022 (.Y (nx6021), .A0 (nx6405), .A1 (nx8158), .B0 (nx8142), .B1 (
          nx8150)) ;
    nand02_2x ix8143 (.Y (nx8142), .A0 (nx6017), .A1 (nx6011)) ;
    nor02_2x ix8145 (.Y (nx8144), .A0 (nx6011), .A1 (nx6017)) ;
    aoi21 ix6034 (.Y (nx6033), .A0 (nx6407), .A1 (nx8184), .B0 (nx8178)) ;
    xnor2 ix8185 (.Y (nx8184), .A0 (nx5811), .A1 (nx7980)) ;
    nor03 ix8179 (.Y (nx8178), .A0 (nx6039), .A1 (nx6407), .A2 (nx6415)) ;
    nor02ii ix6040 (.Y (nx6039), .A0 (nx8144), .A1 (nx6041)) ;
    xnor2 ix6042 (.Y (nx6041), .A0 (nx5815), .A1 (nx5819)) ;
    nor02ii ix8171 (.Y (nx8170), .A0 (nx6041), .A1 (nx8144)) ;
    oai22 ix8215 (.Y (nx8214), .A0 (nx6433), .A1 (nx6049), .B0 (nx6051), .B1 (
          nx6053)) ;
    xnor2 ix6050 (.Y (nx6049), .A0 (nx7950), .A1 (nx6395)) ;
    nor02_2x ix6052 (.Y (nx6051), .A0 (nx6415), .A1 (nx8184)) ;
    nand02_2x ix6054 (.Y (nx6053), .A0 (nx6433), .A1 (nx6055)) ;
    nand02_2x ix6056 (.Y (nx6055), .A0 (nx8184), .A1 (nx6415)) ;
    aoi22 ix6060 (.Y (nx6059), .A0 (nx6407), .A1 (nx8236), .B0 (nx8220), .B1 (
          nx8228)) ;
    nand02_2x ix8221 (.Y (nx8220), .A0 (nx6055), .A1 (nx6049)) ;
    nor02_2x ix8223 (.Y (nx8222), .A0 (nx6049), .A1 (nx6055)) ;
    aoi21 ix6072 (.Y (nx6071), .A0 (nx6407), .A1 (nx8262), .B0 (nx8256)) ;
    xnor2 ix8263 (.Y (nx8262), .A0 (nx5797), .A1 (nx7986)) ;
    nor03 ix8257 (.Y (nx8256), .A0 (nx6077), .A1 (nx6407), .A2 (nx6417)) ;
    nor02ii ix6078 (.Y (nx6077), .A0 (nx8222), .A1 (nx6079)) ;
    xnor2 ix6080 (.Y (nx6079), .A0 (nx5801), .A1 (nx5805)) ;
    nor02ii ix8249 (.Y (nx8248), .A0 (nx6079), .A1 (nx8222)) ;
    oai22 ix8293 (.Y (nx8292), .A0 (nx6433), .A1 (nx6087), .B0 (nx6089), .B1 (
          nx6091)) ;
    xnor2 ix6088 (.Y (nx6087), .A0 (nx7944), .A1 (nx6397)) ;
    nor02_2x ix6090 (.Y (nx6089), .A0 (nx6417), .A1 (nx8262)) ;
    nand02_2x ix6092 (.Y (nx6091), .A0 (nx6433), .A1 (nx6093)) ;
    nand02_2x ix6094 (.Y (nx6093), .A0 (nx8262), .A1 (nx6417)) ;
    aoi22 ix6098 (.Y (nx6097), .A0 (nx6409), .A1 (nx8314), .B0 (nx8298), .B1 (
          nx8306)) ;
    nand02_2x ix8299 (.Y (nx8298), .A0 (nx6093), .A1 (nx6087)) ;
    nor02_2x ix8301 (.Y (nx8300), .A0 (nx6087), .A1 (nx6093)) ;
    aoi21 ix6110 (.Y (nx6109), .A0 (nx6409), .A1 (nx8340), .B0 (nx8334)) ;
    xnor2 ix8341 (.Y (nx8340), .A0 (nx5783), .A1 (nx7992)) ;
    nor03 ix8335 (.Y (nx8334), .A0 (nx6115), .A1 (nx6409), .A2 (nx6419)) ;
    nor02ii ix6116 (.Y (nx6115), .A0 (nx8300), .A1 (nx6117)) ;
    xnor2 ix6118 (.Y (nx6117), .A0 (nx5787), .A1 (nx5791)) ;
    nor02ii ix8327 (.Y (nx8326), .A0 (nx6117), .A1 (nx8300)) ;
    oai22 ix8371 (.Y (nx8370), .A0 (nx6435), .A1 (nx6125), .B0 (nx6127), .B1 (
          nx6129)) ;
    xnor2 ix6126 (.Y (nx6125), .A0 (nx7938), .A1 (nx6399)) ;
    nor02_2x ix6128 (.Y (nx6127), .A0 (nx6419), .A1 (nx8340)) ;
    nand02_2x ix6130 (.Y (nx6129), .A0 (nx6435), .A1 (nx6131)) ;
    nand02_2x ix6132 (.Y (nx6131), .A0 (nx8340), .A1 (nx6419)) ;
    aoi22 ix6136 (.Y (nx6135), .A0 (nx6409), .A1 (nx8392), .B0 (nx8376), .B1 (
          nx8384)) ;
    nand02_2x ix8377 (.Y (nx8376), .A0 (nx6131), .A1 (nx6125)) ;
    nor02_2x ix8379 (.Y (nx8378), .A0 (nx6125), .A1 (nx6131)) ;
    aoi21 ix6148 (.Y (nx6147), .A0 (nx6409), .A1 (nx8418), .B0 (nx8412)) ;
    xnor2 ix8419 (.Y (nx8418), .A0 (nx5769), .A1 (nx7998)) ;
    nor03 ix8413 (.Y (nx8412), .A0 (nx6153), .A1 (nx6411), .A2 (nx6421)) ;
    nor02ii ix6154 (.Y (nx6153), .A0 (nx8378), .A1 (nx6155)) ;
    xnor2 ix6156 (.Y (nx6155), .A0 (nx5773), .A1 (nx5777)) ;
    nor02ii ix8405 (.Y (nx8404), .A0 (nx6155), .A1 (nx8378)) ;
    oai22 ix8449 (.Y (nx8448), .A0 (nx6435), .A1 (nx6163), .B0 (nx6165), .B1 (
          nx6167)) ;
    xnor2 ix6164 (.Y (nx6163), .A0 (nx7932), .A1 (nx6401)) ;
    nor02_2x ix6166 (.Y (nx6165), .A0 (nx6421), .A1 (nx8418)) ;
    nand02_2x ix6168 (.Y (nx6167), .A0 (nx6435), .A1 (nx6169)) ;
    nand02_2x ix6170 (.Y (nx6169), .A0 (nx8418), .A1 (nx6421)) ;
    aoi22 ix6174 (.Y (nx6173), .A0 (nx6411), .A1 (nx8470), .B0 (nx8454), .B1 (
          nx8462)) ;
    nand02_2x ix8455 (.Y (nx8454), .A0 (nx6169), .A1 (nx6163)) ;
    nor02_2x ix8457 (.Y (nx8456), .A0 (nx6163), .A1 (nx6169)) ;
    aoi21 ix6186 (.Y (nx6185), .A0 (nx6411), .A1 (nx8496), .B0 (nx8490)) ;
    xnor2 ix8497 (.Y (nx8496), .A0 (nx5755), .A1 (nx8004)) ;
    nor03 ix8491 (.Y (nx8490), .A0 (nx6191), .A1 (nx6411), .A2 (nx6423)) ;
    nor02ii ix6192 (.Y (nx6191), .A0 (nx8456), .A1 (nx6193)) ;
    xnor2 ix6194 (.Y (nx6193), .A0 (nx5759), .A1 (nx5763)) ;
    nor02ii ix8483 (.Y (nx8482), .A0 (nx6193), .A1 (nx8456)) ;
    oai22 ix8527 (.Y (nx8526), .A0 (nx6435), .A1 (nx6201), .B0 (nx6203), .B1 (
          nx6205)) ;
    xnor2 ix6202 (.Y (nx6201), .A0 (nx7926), .A1 (nx6403)) ;
    nor02_2x ix6204 (.Y (nx6203), .A0 (nx6423), .A1 (nx8496)) ;
    nand02_2x ix6206 (.Y (nx6205), .A0 (nx6435), .A1 (nx6207)) ;
    nand02_2x ix6208 (.Y (nx6207), .A0 (nx8496), .A1 (nx6423)) ;
    aoi22 ix6212 (.Y (nx6211), .A0 (nx6411), .A1 (nx8548), .B0 (nx8532), .B1 (
          nx8540)) ;
    nand02_2x ix8533 (.Y (nx8532), .A0 (nx6207), .A1 (nx6201)) ;
    nor02_2x ix8535 (.Y (nx8534), .A0 (nx6201), .A1 (nx6207)) ;
    aoi21 ix6224 (.Y (nx6223), .A0 (nx6481), .A1 (nx8574), .B0 (nx8568)) ;
    xnor2 ix8575 (.Y (nx8574), .A0 (nx5741), .A1 (nx8010)) ;
    nor03 ix8569 (.Y (nx8568), .A0 (nx6229), .A1 (nx6481), .A2 (nx6425)) ;
    nor02ii ix6230 (.Y (nx6229), .A0 (nx8534), .A1 (nx6231)) ;
    xnor2 ix6232 (.Y (nx6231), .A0 (nx5745), .A1 (nx5749)) ;
    nor02ii ix8561 (.Y (nx8560), .A0 (nx6231), .A1 (nx8534)) ;
    oai22 ix8599 (.Y (nx8598), .A0 (nx6239), .A1 (nx6241), .B0 (nx6481), .B1 (
          nx6243)) ;
    nor02_2x ix6240 (.Y (nx6239), .A0 (nx8012), .A1 (nx7920)) ;
    nand02_2x ix6242 (.Y (nx6241), .A0 (nx5735), .A1 (nx6481)) ;
    xnor2 ix6244 (.Y (nx6243), .A0 (nx8574), .A1 (nx6425)) ;
    aoi32 ix6248 (.Y (nx6247), .A0 (nx8614), .A1 (nx6251), .A2 (nx8776), .B0 (
          overflow), .B1 (nx6257)) ;
    nand02_2x ix6252 (.Y (nx6251), .A0 (nx6481), .A1 (nx1329)) ;
    nand03 ix6256 (.Y (nx6255), .A0 (nx1245), .A1 (input_a[30]), .A2 (
           input_b[30])) ;
    aoi32 ix6262 (.Y (nx6261), .A0 (nx8794), .A1 (nx6267), .A2 (nx8776), .B0 (
          overflow), .B1 (nx6257)) ;
    nand02_2x ix8795 (.Y (nx8794), .A0 (nx6251), .A1 (nx6265)) ;
    xnor2 ix6266 (.Y (nx6265), .A0 (nx1329), .A1 (nx1333)) ;
    aoi32 ix6272 (.Y (nx6271), .A0 (nx8812), .A1 (nx1323), .A2 (nx8776), .B0 (
          overflow), .B1 (nx6257)) ;
    or02 ix8813 (.Y (nx8812), .A0 (nx8746), .A1 (nx8738)) ;
    oai32 ix8843 (.Y (nx8842), .A0 (nx6279), .A1 (nx6429), .A2 (nx6453), .B0 (
          nx6255), .B1 (nx6314)) ;
    nor02ii ix6280 (.Y (nx6279), .A0 (nx8732), .A1 (nx1323)) ;
    aoi32 ix6286 (.Y (nx6285), .A0 (nx8848), .A1 (nx1317), .A2 (nx8776), .B0 (
          overflow), .B1 (nx6257)) ;
    or02 ix8849 (.Y (nx8848), .A0 (nx6429), .A1 (nx8726)) ;
    oai32 ix8879 (.Y (nx8878), .A0 (nx6293), .A1 (nx6431), .A2 (nx6453), .B0 (
          nx6255), .B1 (nx6314)) ;
    nor02ii ix6294 (.Y (nx6293), .A0 (nx8720), .A1 (nx1317)) ;
    aoi32 ix6298 (.Y (nx6297), .A0 (nx8884), .A1 (nx1311), .A2 (nx8776), .B0 (
          overflow), .B1 (nx6257)) ;
    or02 ix8885 (.Y (nx8884), .A0 (nx6431), .A1 (nx8714)) ;
    ao21 ix6304 (.Y (nx6303), .A0 (nx6255), .A1 (nx1245), .B0 (nx6314)) ;
    xnor2 ix6308 (.Y (nx6307), .A0 (input_a[31]), .A1 (input_b[31])) ;
    inv02 ix6268 (.Y (nx6267), .A (nx8746)) ;
    inv02 ix8621 (.Y (nx8620), .A (nx1301)) ;
    inv02 ix8611 (.Y (nx8610), .A (nx1329)) ;
    inv02 ix8605 (.Y (nx8604), .A (nx1331)) ;
    inv02 ix8549 (.Y (nx8548), .A (nx6231)) ;
    inv02 ix8471 (.Y (nx8470), .A (nx6193)) ;
    inv02 ix8393 (.Y (nx8392), .A (nx6155)) ;
    inv02 ix8315 (.Y (nx8314), .A (nx6117)) ;
    inv02 ix8237 (.Y (nx8236), .A (nx6079)) ;
    inv02 ix8159 (.Y (nx8158), .A (nx6041)) ;
    inv02 ix8081 (.Y (nx8080), .A (nx6003)) ;
    inv02 ix8055 (.Y (nx8054), .A (nx5989)) ;
    inv02 ix8017 (.Y (nx8016), .A (nx1341)) ;
    inv02 ix7905 (.Y (nx7904), .A (nx5747)) ;
    inv02 ix2264 (.Y (nx2263), .A (nx7892)) ;
    inv02 ix7881 (.Y (nx7880), .A (nx5775)) ;
    inv02 ix3344 (.Y (nx3343), .A (nx7868)) ;
    inv02 ix7857 (.Y (nx7856), .A (nx5803)) ;
    inv02 ix4424 (.Y (nx4423), .A (nx7844)) ;
    inv02 ix7833 (.Y (nx7832), .A (nx5831)) ;
    inv02 ix5518 (.Y (nx5517), .A (nx7794)) ;
    inv02 ix5532 (.Y (nx5531), .A (nx7750)) ;
    inv02 ix5538 (.Y (nx5537), .A (nx7696)) ;
    inv02 ix7693 (.Y (nx7692), .A (nx5539)) ;
    inv02 ix5554 (.Y (nx5553), .A (nx7624)) ;
    inv02 ix5560 (.Y (nx5559), .A (nx7542)) ;
    inv02 ix5574 (.Y (nx5573), .A (nx7442)) ;
    inv02 ix5562 (.Y (nx5561), .A (nx7440)) ;
    inv02 ix5582 (.Y (nx5581), .A (nx7332)) ;
    inv02 ix5596 (.Y (nx5595), .A (nx7204)) ;
    inv02 ix5602 (.Y (nx5601), .A (nx7066)) ;
    inv02 ix7063 (.Y (nx7062), .A (nx5603)) ;
    inv02 ix5618 (.Y (nx5617), .A (nx6910)) ;
    inv02 ix5624 (.Y (nx5623), .A (nx6744)) ;
    inv02 ix5638 (.Y (nx5637), .A (nx6560)) ;
    inv02 ix5626 (.Y (nx5625), .A (nx6558)) ;
    inv02 ix5646 (.Y (nx5645), .A (nx6366)) ;
    inv02 ix5660 (.Y (nx5659), .A (nx6154)) ;
    inv02 ix5666 (.Y (nx5665), .A (nx5932)) ;
    inv02 ix5929 (.Y (nx5928), .A (nx5667)) ;
    inv02 ix5682 (.Y (nx5681), .A (nx5692)) ;
    inv02 ix5688 (.Y (nx5687), .A (nx5442)) ;
    inv02 ix5702 (.Y (nx5701), .A (nx5174)) ;
    inv02 ix5690 (.Y (nx5689), .A (nx5172)) ;
    inv02 ix5710 (.Y (nx5709), .A (nx4896)) ;
    inv02 ix5724 (.Y (nx5723), .A (nx4600)) ;
    inv02 ix5730 (.Y (nx5729), .A (nx4294)) ;
    inv02 ix4291 (.Y (nx4290), .A (nx5731)) ;
    inv02 ix5148 (.Y (nx5147), .A (nx3920)) ;
    inv02 ix3797 (.Y (nx3796), .A (nx1617)) ;
    inv02 ix8765 (.Y (overflow), .A (nx6255)) ;
    inv02 ix6258 (.Y (nx6257), .A (underflow)) ;
    inv02 ix6313 (.Y (nx6314), .A (nx6257)) ;
    inv02 ix6315 (.Y (nx6316), .A (nx252)) ;
    buf02 ix6370 (.Y (nx6371), .A (nx4202)) ;
    buf02 ix6372 (.Y (nx6373), .A (nx4210)) ;
    buf02 ix6374 (.Y (nx6375), .A (nx4218)) ;
    buf02 ix6376 (.Y (nx6377), .A (nx4226)) ;
    buf02 ix6378 (.Y (nx6379), .A (nx4234)) ;
    buf02 ix6380 (.Y (nx6381), .A (nx4242)) ;
    buf02 ix6382 (.Y (nx6383), .A (nx4250)) ;
    buf02 ix6384 (.Y (nx6385), .A (nx4258)) ;
    buf02 ix6386 (.Y (nx6387), .A (nx4266)) ;
    buf02 ix6388 (.Y (nx6389), .A (nx4274)) ;
    buf02 ix6390 (.Y (nx6391), .A (nx7970)) ;
    buf02 ix6392 (.Y (nx6393), .A (nx7976)) ;
    buf02 ix6394 (.Y (nx6395), .A (nx7982)) ;
    buf02 ix6396 (.Y (nx6397), .A (nx7988)) ;
    buf02 ix6398 (.Y (nx6399), .A (nx7994)) ;
    buf02 ix6400 (.Y (nx6401), .A (nx8000)) ;
    buf02 ix6402 (.Y (nx6403), .A (nx8006)) ;
    inv02 ix6404 (.Y (nx6405), .A (nx6491)) ;
    inv02 ix6406 (.Y (nx6407), .A (nx6491)) ;
    inv02 ix6408 (.Y (nx6409), .A (nx6491)) ;
    inv02 ix6410 (.Y (nx6411), .A (nx6491)) ;
    buf02 ix6412 (.Y (nx6413), .A (nx8092)) ;
    buf02 ix6414 (.Y (nx6415), .A (nx8170)) ;
    buf02 ix6416 (.Y (nx6417), .A (nx8248)) ;
    buf02 ix6418 (.Y (nx6419), .A (nx8326)) ;
    buf02 ix6420 (.Y (nx6421), .A (nx8404)) ;
    buf02 ix6422 (.Y (nx6423), .A (nx8482)) ;
    buf02 ix6424 (.Y (nx6425), .A (nx8560)) ;
    buf02 ix6426 (.Y (nx6427), .A (nx8638)) ;
    buf02 ix6428 (.Y (nx6429), .A (nx8750)) ;
    buf02 ix6430 (.Y (nx6431), .A (nx8754)) ;
    inv02 ix6432 (.Y (nx6433), .A (nx6481)) ;
    inv02 ix6434 (.Y (nx6435), .A (nx6481)) ;
    inv02 ix6436 (.Y (nx6437), .A (nx8016)) ;
    inv02 ix6440 (.Y (nx6441), .A (input_a[1])) ;
    inv02 ix6446 (.Y (nx6447), .A (input_a[0])) ;
    inv02 ix6452 (.Y (nx6453), .A (nx8776)) ;
    ao32 ix4275 (.Y (nx4274), .A0 (input_b[22]), .A1 (input_a[21]), .A2 (
         input_a[20]), .B0 (nx6460), .B1 (nx4038)) ;
    inv02 ix6459 (.Y (nx6460), .A (nx1359)) ;
    ao32 ix4267 (.Y (nx4266), .A0 (input_b[22]), .A1 (input_a[19]), .A2 (
         input_a[18]), .B0 (nx6462), .B1 (nx4054)) ;
    inv02 ix6461 (.Y (nx6462), .A (nx1367)) ;
    ao32 ix4259 (.Y (nx4258), .A0 (input_b[22]), .A1 (input_a[17]), .A2 (
         input_a[16]), .B0 (nx6464), .B1 (nx4070)) ;
    inv02 ix6463 (.Y (nx6464), .A (nx1375)) ;
    ao32 ix4251 (.Y (nx4250), .A0 (input_b[22]), .A1 (input_a[15]), .A2 (
         input_a[14]), .B0 (nx6466), .B1 (nx4086)) ;
    inv02 ix6465 (.Y (nx6466), .A (nx1383)) ;
    ao32 ix4243 (.Y (nx4242), .A0 (input_b[22]), .A1 (input_a[13]), .A2 (
         input_a[12]), .B0 (nx6468), .B1 (nx4102)) ;
    inv02 ix6467 (.Y (nx6468), .A (nx1391)) ;
    ao32 ix4235 (.Y (nx4234), .A0 (input_b[22]), .A1 (input_a[11]), .A2 (
         input_a[10]), .B0 (nx6470), .B1 (nx4118)) ;
    inv02 ix6469 (.Y (nx6470), .A (nx1399)) ;
    ao32 ix4227 (.Y (nx4226), .A0 (input_b[22]), .A1 (input_a[9]), .A2 (
         input_a[8]), .B0 (nx6472), .B1 (nx4134)) ;
    inv02 ix6471 (.Y (nx6472), .A (nx1407)) ;
    ao32 ix4219 (.Y (nx4218), .A0 (input_b[22]), .A1 (input_a[7]), .A2 (
         input_a[6]), .B0 (nx6475), .B1 (nx4150)) ;
    inv02 ix6473 (.Y (nx6475), .A (nx1415)) ;
    ao32 ix4211 (.Y (nx4210), .A0 (input_b[22]), .A1 (input_a[5]), .A2 (
         input_a[4]), .B0 (nx6477), .B1 (nx4166)) ;
    inv02 ix6476 (.Y (nx6477), .A (nx1423)) ;
    ao32 ix4203 (.Y (nx4202), .A0 (input_b[22]), .A1 (input_a[3]), .A2 (
         input_a[2]), .B0 (nx6479), .B1 (nx4182)) ;
    inv02 ix6478 (.Y (nx6479), .A (nx1431)) ;
    and03 ix3191 (.Y (nx3190), .A0 (input_a[1]), .A1 (input_b[22]), .A2 (
          input_a[0])) ;
    and04 ix3193 (.Y (nx3192), .A0 (input_b[21]), .A1 (input_a[1]), .A2 (
          input_b[22]), .A3 (input_a[0])) ;
    nor02ii ix2171 (.Y (nx2170), .A0 (nx1985), .A1 (nx2009)) ;
    nand04 ix2161 (.Y (nx2009), .A0 (input_b[19]), .A1 (input_b[20]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix1992 (.Y (nx1991), .A0 (nx2009), .A1 (nx2662)) ;
    nor02ii ix2659 (.Y (nx2658), .A0 (nx1999), .A1 (nx1589)) ;
    nand04 ix2649 (.Y (nx1589), .A0 (input_b[20]), .A1 (input_b[21]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix3209 (.Y (nx3208), .A0 (nx1589), .A1 (nx1593)) ;
    nor02ii ix1363 (.Y (nx1362), .A0 (nx2343), .A1 (nx2369)) ;
    nand04 ix1353 (.Y (nx2369), .A0 (input_b[17]), .A1 (input_b[18]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix2350 (.Y (nx2349), .A0 (nx2369), .A1 (nx1742)) ;
    nor02ii ix1739 (.Y (nx1738), .A0 (nx2357), .A1 (nx1973)) ;
    nand04 ix1729 (.Y (nx1973), .A0 (input_b[18]), .A1 (input_b[19]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix2374 (.Y (nx2373), .A0 (nx1973), .A1 (nx2174)) ;
    nor02ii ix779 (.Y (nx778), .A0 (nx2701), .A1 (nx2727)) ;
    nand04 ix769 (.Y (nx2727), .A0 (input_b[15]), .A1 (input_b[16]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix2708 (.Y (nx2707), .A0 (nx2727), .A1 (nx1046)) ;
    nor02ii ix1043 (.Y (nx1042), .A0 (nx2715), .A1 (nx2331)) ;
    nand04 ix1033 (.Y (nx2331), .A0 (input_b[16]), .A1 (input_b[17]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix2732 (.Y (nx2731), .A0 (nx2331), .A1 (nx1366)) ;
    nor02ii ix419 (.Y (nx418), .A0 (nx3059), .A1 (nx3085)) ;
    nand04 ix409 (.Y (nx3085), .A0 (input_b[13]), .A1 (input_b[14]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix3066 (.Y (nx3065), .A0 (nx3085), .A1 (nx574)) ;
    nor02ii ix571 (.Y (nx570), .A0 (nx3073), .A1 (nx2689)) ;
    nand04 ix561 (.Y (nx2689), .A0 (input_b[14]), .A1 (input_b[15]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix3090 (.Y (nx3089), .A0 (nx2689), .A1 (nx782)) ;
    nor02ii ix291 (.Y (nx290), .A0 (nx3417), .A1 (nx3443)) ;
    nand04 ix281 (.Y (nx3443), .A0 (input_b[11]), .A1 (input_b[12]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix3424 (.Y (nx3423), .A0 (nx3443), .A1 (nx326)) ;
    nor02ii ix323 (.Y (nx322), .A0 (nx3431), .A1 (nx3047)) ;
    nand04 ix313 (.Y (nx3047), .A0 (input_b[12]), .A1 (input_b[13]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix3448 (.Y (nx3447), .A0 (nx3047), .A1 (nx422)) ;
    nor02ii ix491 (.Y (nx490), .A0 (nx3775), .A1 (nx3801)) ;
    nand04 ix375 (.Y (nx3801), .A0 (input_b[9]), .A1 (input_b[10]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix3782 (.Y (nx3781), .A0 (nx3801), .A1 (nx364)) ;
    nor02ii ix363 (.Y (nx362), .A0 (nx3789), .A1 (nx3405)) ;
    nand04 ix303 (.Y (nx3405), .A0 (input_b[10]), .A1 (input_b[11]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix3806 (.Y (nx3805), .A0 (nx3405), .A1 (nx292)) ;
    nor02ii ix915 (.Y (nx914), .A0 (nx4133), .A1 (nx4159)) ;
    nand04 ix687 (.Y (nx4159), .A0 (input_b[7]), .A1 (input_b[8]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix4140 (.Y (nx4139), .A0 (nx4159), .A1 (nx676)) ;
    nor02ii ix675 (.Y (nx674), .A0 (nx4147), .A1 (nx3763)) ;
    nand04 ix503 (.Y (nx3763), .A0 (input_b[8]), .A1 (input_b[9]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix4164 (.Y (nx4163), .A0 (nx3763), .A1 (nx492)) ;
    nor02ii ix1563 (.Y (nx1562), .A0 (nx4491), .A1 (nx4517)) ;
    nand04 ix1223 (.Y (nx4517), .A0 (input_b[5]), .A1 (input_b[6]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix4498 (.Y (nx4497), .A0 (nx4517), .A1 (nx1212)) ;
    nor02ii ix1211 (.Y (nx1210), .A0 (nx4505), .A1 (nx4121)) ;
    nand04 ix927 (.Y (nx4121), .A0 (input_b[6]), .A1 (input_b[7]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix4522 (.Y (nx4521), .A0 (nx4121), .A1 (nx916)) ;
    nor02ii ix2435 (.Y (nx2434), .A0 (nx4849), .A1 (nx4875)) ;
    nand04 ix1983 (.Y (nx4875), .A0 (input_b[3]), .A1 (input_b[4]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix4856 (.Y (nx4855), .A0 (nx4875), .A1 (nx1972)) ;
    nor02ii ix1971 (.Y (nx1970), .A0 (nx4863), .A1 (nx4479)) ;
    nand04 ix1575 (.Y (nx4479), .A0 (input_b[4]), .A1 (input_b[5]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix4880 (.Y (nx4879), .A0 (nx4479), .A1 (nx1564)) ;
    nor02ii ix2955 (.Y (nx2954), .A0 (nx5203), .A1 (nx4837)) ;
    nand04 ix2447 (.Y (nx4837), .A0 (input_b[2]), .A1 (input_b[3]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix5210 (.Y (nx5209), .A0 (nx4837), .A1 (nx2436)) ;
    nor02ii ix3531 (.Y (nx3530), .A0 (nx5381), .A1 (nx5193)) ;
    nand04 ix2967 (.Y (nx5193), .A0 (input_b[1]), .A1 (input_b[2]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    xor2 ix5388 (.Y (nx5387), .A0 (nx5193), .A1 (nx2956)) ;
    xor2 ix5906 (.Y (nx5905), .A0 (nx5371), .A1 (nx3532)) ;
    nand04 ix3543 (.Y (nx5371), .A0 (input_b[0]), .A1 (input_b[1]), .A2 (
           input_a[0]), .A3 (input_a[1])) ;
    nor02ii ix8037 (.Y (product[0]), .A0 (nx5959), .A1 (nx6483)) ;
    mux21 ix5960 (.Y (nx5959), .A0 (nx5963), .A1 (nx8028), .S0 (nx8016)) ;
    nor02ii ix8063 (.Y (product[1]), .A0 (nx5967), .A1 (nx6483)) ;
    nor02ii ix8089 (.Y (product[2]), .A0 (nx5981), .A1 (nx6483)) ;
    nor02ii ix8115 (.Y (product[3]), .A0 (nx5995), .A1 (nx6483)) ;
    and02 ix8141 (.Y (product[4]), .A0 (nx6483), .A1 (nx8136)) ;
    nor02ii ix8167 (.Y (product[5]), .A0 (nx6021), .A1 (nx6483)) ;
    nor02ii ix8151 (.Y (nx8150), .A0 (nx8144), .A1 (nx6491)) ;
    nor02ii ix8193 (.Y (product[6]), .A0 (nx6033), .A1 (nx6483)) ;
    and02 ix8219 (.Y (product[7]), .A0 (nx6485), .A1 (nx8214)) ;
    nor02ii ix8245 (.Y (product[8]), .A0 (nx6059), .A1 (nx6485)) ;
    nor02ii ix8229 (.Y (nx8228), .A0 (nx8222), .A1 (nx6491)) ;
    nor02ii ix8271 (.Y (product[9]), .A0 (nx6071), .A1 (nx6485)) ;
    and02 ix8297 (.Y (product[10]), .A0 (nx6485), .A1 (nx8292)) ;
    nor02ii ix8323 (.Y (product[11]), .A0 (nx6097), .A1 (nx6485)) ;
    nor02ii ix8307 (.Y (nx8306), .A0 (nx8300), .A1 (nx6437)) ;
    nor02ii ix8349 (.Y (product[12]), .A0 (nx6109), .A1 (nx6485)) ;
    and02 ix8375 (.Y (product[13]), .A0 (nx6485), .A1 (nx8370)) ;
    nor02ii ix8401 (.Y (product[14]), .A0 (nx6135), .A1 (nx6487)) ;
    nor02ii ix8385 (.Y (nx8384), .A0 (nx8378), .A1 (nx6437)) ;
    nor02ii ix8427 (.Y (product[15]), .A0 (nx6147), .A1 (nx6487)) ;
    and02 ix8453 (.Y (product[16]), .A0 (nx6487), .A1 (nx8448)) ;
    nor02ii ix8479 (.Y (product[17]), .A0 (nx6173), .A1 (nx6487)) ;
    nor02ii ix8463 (.Y (nx8462), .A0 (nx8456), .A1 (nx6437)) ;
    nor02ii ix8505 (.Y (product[18]), .A0 (nx6185), .A1 (nx6487)) ;
    and02 ix8531 (.Y (product[19]), .A0 (nx6487), .A1 (nx8526)) ;
    nor02ii ix8557 (.Y (product[20]), .A0 (nx6211), .A1 (nx6487)) ;
    nor02ii ix8541 (.Y (nx8540), .A0 (nx8534), .A1 (nx6437)) ;
    nor02ii ix8583 (.Y (product[21]), .A0 (nx6223), .A1 (nx6489)) ;
    and02 ix8603 (.Y (product[22]), .A0 (nx6489), .A1 (nx8598)) ;
    nor02ii ix8793 (.Y (product[23]), .A0 (nx6247), .A1 (nx6489)) ;
    or02 ix8615 (.Y (nx8614), .A0 (nx1329), .A1 (nx8016)) ;
    nor02ii ix8811 (.Y (product[24]), .A0 (nx6261), .A1 (nx6489)) ;
    nor02ii ix8829 (.Y (product[25]), .A0 (nx6271), .A1 (nx6489)) ;
    and02 ix8847 (.Y (product[26]), .A0 (nx6489), .A1 (nx8842)) ;
    nand02_2x ix6282 (.Y (nx8776), .A0 (nx6255), .A1 (nx6314)) ;
    nor02ii ix8865 (.Y (product[27]), .A0 (nx6285), .A1 (nx6489)) ;
    and02 ix8883 (.Y (product[28]), .A0 (nx6316), .A1 (nx8878)) ;
    nor02ii ix8901 (.Y (product[29]), .A0 (nx6297), .A1 (nx6316)) ;
    nor02ii ix8913 (.Y (product[30]), .A0 (nx6303), .A1 (nx6316)) ;
    nor02ii ix8919 (.Y (product[31]), .A0 (nx6307), .A1 (nx6316)) ;
    inv02 ix6480 (.Y (nx6481), .A (nx1341)) ;
    inv02 ix6482 (.Y (nx6483), .A (nx252)) ;
    inv02 ix6484 (.Y (nx6485), .A (nx252)) ;
    inv02 ix6486 (.Y (nx6487), .A (nx252)) ;
    inv02 ix6488 (.Y (nx6489), .A (nx252)) ;
    inv02 ix6490 (.Y (nx6491), .A (nx8016)) ;
endmodule

